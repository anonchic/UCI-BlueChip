-- DDR controller
  constant CFG_DDR2SP  		       : integer := CONFIG_DDR2SP;
  constant CFG_DDR2SP_INIT  	   : integer := CONFIG_DDR2SP_INIT;
  constant CFG_DDR2SP_FREQ   	   : integer := CONFIG_DDR2SP_FREQ;
  constant CFG_DDR2SP_DATAWIDTH  : integer := CONFIG_DDR2SP_DATAWIDTH;
  constant CFG_DDR2SP_COL    	   : integer := CONFIG_DDR2SP_COL;
  constant CFG_DDR2SP_SIZE  	   : integer := CONFIG_DDR2SP_MBYTE;
  constant CFG_DDR2SP_DELAY0 	   : integer := CONFIG_DDR2SP_DELAY0;
  constant CFG_DDR2SP_DELAY1 	   : integer := CONFIG_DDR2SP_DELAY1;
  constant CFG_DDR2SP_DELAY2 	   : integer := CONFIG_DDR2SP_DELAY2;
  constant CFG_DDR2SP_DELAY3 	   : integer := CONFIG_DDR2SP_DELAY3;
  constant CFG_DDR2SP_DELAY4 	   : integer := CONFIG_DDR2SP_DELAY4;
  constant CFG_DDR2SP_DELAY5 	   : integer := CONFIG_DDR2SP_DELAY5;
  constant CFG_DDR2SP_DELAY6 	   : integer := CONFIG_DDR2SP_DELAY6;
  constant CFG_DDR2SP_DELAY7 	   : integer := CONFIG_DDR2SP_DELAY7;

