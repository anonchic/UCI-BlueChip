package memoryPreLoad is
    CONSTANT NAHBMST : integer := 16;
    CONSTANT NAHBSLV : integer := 16;
    CONSTANT NAPBSLV : integer := 16;
    CONSTANT NAHBIRQ : integer := 32;
    CONSTANT NAHBAMR : integer := 4;
    CONSTANT NAHBIR : integer := 4;
    CONSTANT NAHBCFG : integer := 4 + 4;
    CONSTANT NAPBIR : integer := 1;
    CONSTANT NAPBAMR : integer := 1;
    CONSTANT NAPBCFG : integer := 1 + 1;
    CONSTANT NBUS : integer := 4;
    SUBTYPE amba_config_word IS std_logic_vector ( 31 downto 0 );
    TYPE ahb_config_type IS ARRAY ( 0 to 4 + 4 - 1 ) OF amba_config_word;
    TYPE apb_config_type IS ARRAY ( 0 to 1 + 1 - 1 ) OF amba_config_word;
    TYPE ahb_mst_in_type IS RECORD
        hgrant : std_logic_vector ( 0 to 16 - 1 );
        hready : std_ulogic;
        hresp : std_logic_vector ( 1 downto 0 );
        hrdata : std_logic_vector ( 31 downto 0 );
        hcache : std_ulogic;
        hirq : std_logic_vector ( 32 - 1 downto 0 );
        testen : std_ulogic;
        testrst : std_ulogic;
        scanen : std_ulogic;
        testoen : std_ulogic;
    END RECORD;
    TYPE ahb_mst_out_type IS RECORD
        hbusreq : std_ulogic;
        hlock : std_ulogic;
        htrans : std_logic_vector ( 1 downto 0 );
        haddr : std_logic_vector ( 31 downto 0 );
        hwrite : std_ulogic;
        hsize : std_logic_vector ( 2 downto 0 );
        hburst : std_logic_vector ( 2 downto 0 );
        hprot : std_logic_vector ( 3 downto 0 );
        hwdata : std_logic_vector ( 31 downto 0 );
        hirq : std_logic_vector ( 32 - 1 downto 0 );
        hconfig : ahb_config_type;
        hindex : integer RANGE 0 to 16 - 1;
    END RECORD;
    TYPE ahb_slv_in_type IS RECORD
        hsel : std_logic_vector ( 0 to 16 - 1 );
        haddr : std_logic_vector ( 31 downto 0 );
        hwrite : std_ulogic;
        htrans : std_logic_vector ( 1 downto 0 );
        hsize : std_logic_vector ( 2 downto 0 );
        hburst : std_logic_vector ( 2 downto 0 );
        hwdata : std_logic_vector ( 31 downto 0 );
        hprot : std_logic_vector ( 3 downto 0 );
        hready : std_ulogic;
        hmaster : std_logic_vector ( 3 downto 0 );
        hmastlock : std_ulogic;
        hmbsel : std_logic_vector ( 0 to 4 - 1 );
        hcache : std_ulogic;
        hirq : std_logic_vector ( 32 - 1 downto 0 );
        testen : std_ulogic;
        testrst : std_ulogic;
        scanen : std_ulogic;
        testoen : std_ulogic;
    END RECORD;
    TYPE ahb_slv_out_type IS RECORD
        hready : std_ulogic;
        hresp : std_logic_vector ( 1 downto 0 );
        hrdata : std_logic_vector ( 31 downto 0 );
        hsplit : std_logic_vector ( 15 downto 0 );
        hcache : std_ulogic;
        hirq : std_logic_vector ( 32 - 1 downto 0 );
        hconfig : ahb_config_type;
        hindex : integer RANGE 0 to 16 - 1;
    END RECORD;
    TYPE ahb_mst_out_vector_type IS ARRAY ( natural RANGE <> ) OF ahb_mst_out_type;
    TYPE ahb_slv_out_vector_type IS ARRAY ( natural RANGE <> ) OF ahb_slv_out_type;
    SUBTYPE ahb_mst_out_vector IS ahb_mst_out_vector_type ( 16 - 1 downto 0 );
    SUBTYPE ahb_slv_out_vector IS ahb_slv_out_vector_type ( 16 - 1 downto 0 );
    TYPE ahb_mst_out_bus_vector IS ARRAY ( 0 to 4 - 1 ) OF ahb_mst_out_vector;
    TYPE ahb_slv_out_bus_vector IS ARRAY ( 0 to 4 - 1 ) OF ahb_slv_out_vector;
    CONSTANT HTRANS_IDLE : std_logic_vector ( 1 downto 0 ) := "00";
    CONSTANT HTRANS_BUSY : std_logic_vector ( 1 downto 0 ) := "01";
    CONSTANT HTRANS_NONSEQ : std_logic_vector ( 1 downto 0 ) := "10";
    CONSTANT HTRANS_SEQ : std_logic_vector ( 1 downto 0 ) := "11";
    CONSTANT HBURST_SINGLE : std_logic_vector ( 2 downto 0 ) := "000";
    CONSTANT HBURST_INCR : std_logic_vector ( 2 downto 0 ) := "001";
    CONSTANT HBURST_WRAP4 : std_logic_vector ( 2 downto 0 ) := "010";
    CONSTANT HBURST_INCR4 : std_logic_vector ( 2 downto 0 ) := "011";
    CONSTANT HBURST_WRAP8 : std_logic_vector ( 2 downto 0 ) := "100";
    CONSTANT HBURST_INCR8 : std_logic_vector ( 2 downto 0 ) := "101";
    CONSTANT HBURST_WRAP16 : std_logic_vector ( 2 downto 0 ) := "110";
    CONSTANT HBURST_INCR16 : std_logic_vector ( 2 downto 0 ) := "111";
    CONSTANT HSIZE_BYTE : std_logic_vector ( 2 downto 0 ) := "000";
    CONSTANT HSIZE_HWORD : std_logic_vector ( 2 downto 0 ) := "001";
    CONSTANT HSIZE_WORD : std_logic_vector ( 2 downto 0 ) := "010";
    CONSTANT HSIZE_DWORD : std_logic_vector ( 2 downto 0 ) := "011";
    CONSTANT HSIZE_4WORD : std_logic_vector ( 2 downto 0 ) := "100";
    CONSTANT HSIZE_8WORD : std_logic_vector ( 2 downto 0 ) := "101";
    CONSTANT HSIZE_16WORD : std_logic_vector ( 2 downto 0 ) := "110";
    CONSTANT HSIZE_32WORD : std_logic_vector ( 2 downto 0 ) := "111";
    CONSTANT HRESP_OKAY : std_logic_vector ( 1 downto 0 ) := "00";
    CONSTANT HRESP_ERROR : std_logic_vector ( 1 downto 0 ) := "01";
    CONSTANT HRESP_RETRY : std_logic_vector ( 1 downto 0 ) := "10";
    CONSTANT HRESP_SPLIT : std_logic_vector ( 1 downto 0 ) := "11";
    TYPE apb_slv_in_type IS RECORD
        psel : std_logic_vector ( 0 to 16 - 1 );
        penable : std_ulogic;
        paddr : std_logic_vector ( 31 downto 0 );
        pwrite : std_ulogic;
        pwdata : std_logic_vector ( 31 downto 0 );
        pirq : std_logic_vector ( 32 - 1 downto 0 );
        testen : std_ulogic;
        testrst : std_ulogic;
        scanen : std_ulogic;
        testoen : std_ulogic;
    END RECORD;
    TYPE apb_slv_out_type IS RECORD
        prdata : std_logic_vector ( 31 downto 0 );
        pirq : std_logic_vector ( 32 - 1 downto 0 );
        pconfig : apb_config_type;
        pindex : integer RANGE 0 to 16 - 1;
    END RECORD;
    TYPE apb_slv_out_vector IS ARRAY ( 0 to 16 - 1 ) OF apb_slv_out_type;
    CONSTANT AMBA_CONFIG_VER0 : std_logic_vector ( 1 downto 0 ) := "00";
    SUBTYPE amba_vendor_type IS integer RANGE 0 to 16#ff#;
    SUBTYPE amba_device_type IS integer RANGE 0 to 16#3ff#;
    SUBTYPE amba_version_type IS integer RANGE 0 to 16#3f#;
    SUBTYPE amba_cfgver_type IS integer RANGE 0 to 3;
    SUBTYPE amba_irq_type IS integer RANGE 0 to 32 - 1;
    SUBTYPE ahb_addr_type IS integer RANGE 0 to 16#fff#;
    CONSTANT zx : std_logic_vector ( 31 downto 0 ) := ( OTHERS => '0' );
    CONSTANT zxirq : std_logic_vector ( 32 - 1 downto 0 ) := ( OTHERS => '0' );
    CONSTANT zy : std_logic_vector ( 0 to 31 ) := ( OTHERS => '0' );
    TYPE memory_in_type IS RECORD
        data : std_logic_vector ( 31 downto 0 );
        brdyn : std_logic;
        bexcn : std_logic;
        writen : std_logic;
        wrn : std_logic_vector ( 3 downto 0 );
        bwidth : std_logic_vector ( 1 downto 0 );
        sd : std_logic_vector ( 63 downto 0 );
        cb : std_logic_vector ( 7 downto 0 );
        scb : std_logic_vector ( 7 downto 0 );
        edac : std_logic;
    END RECORD;
    TYPE memory_out_type IS RECORD
        address : std_logic_vector ( 31 downto 0 );
        data : std_logic_vector ( 31 downto 0 );
        sddata : std_logic_vector ( 63 downto 0 );
        ramsn : std_logic_vector ( 7 downto 0 );
        ramoen : std_logic_vector ( 7 downto 0 );
        ramn : std_ulogic;
        romn : std_ulogic;
        mben : std_logic_vector ( 3 downto 0 );
        iosn : std_logic;
        romsn : std_logic_vector ( 7 downto 0 );
        oen : std_logic;
        writen : std_logic;
        wrn : std_logic_vector ( 3 downto 0 );
        bdrive : std_logic_vector ( 3 downto 0 );
        vbdrive : std_logic_vector ( 31 downto 0 );
        svbdrive : std_logic_vector ( 63 downto 0 );
        read : std_logic;
        sa : std_logic_vector ( 14 downto 0 );
        cb : std_logic_vector ( 7 downto 0 );
        scb : std_logic_vector ( 7 downto 0 );
        vcdrive : std_logic_vector ( 7 downto 0 );
        svcdrive : std_logic_vector ( 7 downto 0 );
        ce : std_ulogic;
    END RECORD;
    TYPE sdctrl_in_type IS RECORD
        wprot : std_ulogic;
        data : std_logic_vector ( 127 downto 0 );
        cb : std_logic_vector ( 15 downto 0 );
    END RECORD;
    TYPE sdctrl_out_type IS RECORD
        sdcke : std_logic_vector ( 1 downto 0 );
        sdcsn : std_logic_vector ( 1 downto 0 );
        sdwen : std_ulogic;
        rasn : std_ulogic;
        casn : std_ulogic;
        dqm : std_logic_vector ( 15 downto 0 );
        bdrive : std_ulogic;
        qdrive : std_ulogic;
        vbdrive : std_logic_vector ( 31 downto 0 );
        address : std_logic_vector ( 16 downto 2 );
        data : std_logic_vector ( 127 downto 0 );
        cb : std_logic_vector ( 15 downto 0 );
        ce : std_ulogic;
        ba : std_logic_vector ( 1 downto 0 );
        cal_en : std_logic_vector ( 7 downto 0 );
        cal_inc : std_logic_vector ( 7 downto 0 );
        cal_rst : std_logic;
        odt : std_logic_vector ( 1 downto 0 );
    END RECORD;
    TYPE sdram_out_type IS RECORD
        sdcke : std_logic_vector ( 1 downto 0 );
        sdcsn : std_logic_vector ( 1 downto 0 );
        sdwen : std_ulogic;
        rasn : std_ulogic;
        casn : std_ulogic;
        dqm : std_logic_vector ( 7 downto 0 );
    END RECORD;
end package memoryPreLoad;
