------------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2003 - 2008, Gaisler Research
--  Copyright (C) 2008, 2009, Aeroflex Gaisler
--
--  This program is free software; you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation; either version 2 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 
-----------------------------------------------------------------------------
-- Entity: 	iu3
-- File:	iu3.vhd
-- Author:	Jiri Gaisler, Edvin Catovic, Gaisler Research
-- Description:	LEON3 7-stage integer pipline
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library grlib;
use grlib.sparc.all;
use grlib.stdlib.all;
library techmap;
use techmap.gencomp.all;
library gaisler;
use gaisler.leon3.all;
use gaisler.libiu.all;
use gaisler.arith.all;
-- pragma translate_off
use grlib.sparc_disas.all;
-- pragma translate_on

entity iu3 is
  generic (
    nwin     : integer range 2 to 32 := 8;
    isets    : integer range 1 to 4 := 2;
    dsets    : integer range 1 to 4 := 2;
    fpu      : integer range 0 to 15 := 0;
    v8       : integer range 0 to 63 := 2;
    cp, mac  : integer range 0 to 1 := 0;
    dsu      : integer range 0 to 1 := 1;
    nwp      : integer range 0 to 4 := 2;
    pclow    : integer range 0 to 2 := 2;
    notag    : integer range 0 to 1 := 0;
    index    : integer range 0 to 15:= 0;
    lddel    : integer range 1 to 2 := 1;
    irfwt    : integer range 0 to 1 := 0;
    disas    : integer range 0 to 2 := 0;
    tbuf     : integer range 0 to 64 := 2;  -- trace buf size in kB (0 - no trace buffer)
    pwd      : integer range 0 to 2 := 0;   -- power-down
    svt      : integer range 0 to 1 := 0;   -- single-vector trapping
    rstaddr  : integer := 16#00000#;        -- reset vector MSB address
    smp      : integer range 0 to 15 := 0;  -- support SMP systems
    fabtech  : integer range 0 to NTECH := 20;
    clk2x    : integer := 0
  );
  port (
    clk   : in  std_ulogic;
    rstn  : in  std_ulogic;
    holdn : in  std_ulogic;
    ici   : buffer icache_in_type;
    ico   : in  icache_out_type;
    dci   : buffer dcache_in_type;
    dco   : in  dcache_out_type;
    rfi   : buffer iregfile_in_type;
    rfo   : in  iregfile_out_type;
    irqi  : in  l3_irq_in_type;
    irqo  : buffer l3_irq_out_type;
    dbgi  : in  l3_debug_in_type;
    dbgo  : buffer l3_debug_out_type;
    muli  : buffer mul32_in_type;
    mulo  : in  mul32_out_type;
    divi  : buffer div32_in_type;
    divo  : in  div32_out_type;
    fpo   : in  fpc_out_type;
    fpi   : buffer fpc_in_type;
    cpo   : in  fpc_out_type;
    cpi   : buffer fpc_in_type;
    tbo   : in  tracebuf_out_type;
    tbi   : buffer tracebuf_in_type;
    sclk   : in  std_ulogic
    );
end;

architecture rtl of iu3 is

  constant ISETMSB : integer := 0;
  constant DSETMSB : integer := 0;
  constant RFBITS : integer range 6 to 10 := 8;
  constant NWINLOG2   : integer range 1 to 5 := 3;
  constant CWPOPT : boolean := true;
  constant CWPMIN : std_logic_vector(2 downto 0) := "000";
  constant CWPMAX : std_logic_vector(2 downto 0) := "111";
  constant FPEN   : boolean := (fpu /= 0);
  constant CPEN   : boolean := false;
  constant MULEN  : boolean := true;
  constant MULTYPE: integer := 0;
  constant DIVEN  : boolean := true;
  constant MACEN  : boolean := false;
  constant MACPIPE: boolean := false;
  constant IMPL   : integer := 15;
  constant VER    : integer := 3;
  constant DBGUNIT : boolean := true;
  constant TRACEBUF   : boolean := true;
  constant TBUFBITS : integer := 7;
  constant PWRD1  : boolean := false; --(pwd = 1) and not (index /= 0);
  constant PWRD2  : boolean := false; --(pwd = 2) or (index /= 0);
  constant RS1OPT : boolean := true;
  constant DYNRST : boolean := false;
  
  subtype word is std_logic_vector(31 downto 0);
  subtype pctype is std_logic_vector(31 downto 2);
  subtype rfatype is std_logic_vector(8-1 downto 0);
  subtype cwptype is std_logic_vector(3-1 downto 0);
  type icdtype is array (0 to 2-1) of word;
  type dcdtype is array (0 to 2-1) of word;

  type dc_in_type is record
    signed, enaddr, read, write, lock , dsuen : std_ulogic;
    size : std_logic_vector(1 downto 0);
    asi  : std_logic_vector(7 downto 0);    
  end record;
  
  type pipeline_ctrl_type is record
    pc    : pctype;
    inst  : word;
    cnt   : std_logic_vector(1 downto 0);
    rd    : rfatype;
    tt    : std_logic_vector(5 downto 0);
    trap  : std_ulogic;
    annul : std_ulogic;
    wreg  : std_ulogic;
    wicc  : std_ulogic;
    wy    : std_ulogic;
    ld    : std_ulogic;
    pv    : std_ulogic;
    rett  : std_ulogic;
  end record;
  
  type fetch_reg_type is record
    pc     : pctype;
    branch : std_ulogic;
  end record;
  
  type decode_reg_type is record
    pc    : pctype;
    inst  : icdtype;
    cwp   : cwptype;
    set   : std_logic_vector(0 downto 0);
    mexc  : std_ulogic;
    cnt   : std_logic_vector(1 downto 0);
    pv    : std_ulogic;
    annul : std_ulogic;
    inull : std_ulogic;
    step  : std_ulogic;        
  end record;
  
  type regacc_reg_type is record
    ctrl  : pipeline_ctrl_type;
    rs1   : std_logic_vector(4 downto 0);
    rfa1, rfa2 : rfatype;
    rsel1, rsel2 : std_logic_vector(2 downto 0);
    rfe1, rfe2 : std_ulogic;
    cwp   : cwptype;
    imm   : word;
    ldcheck1 : std_ulogic;
    ldcheck2 : std_ulogic;
    ldchkra : std_ulogic;
    ldchkex : std_ulogic;
    su : std_ulogic;
    et : std_ulogic;
    wovf : std_ulogic;
    wunf : std_ulogic;
    ticc : std_ulogic;
    jmpl : std_ulogic;
    step  : std_ulogic;            
    mulstart : std_ulogic;            
    divstart : std_ulogic;            
  end record;
  
  type execute_reg_type is record
    ctrl   : pipeline_ctrl_type;
    op1    : word;
    op2    : word;
    aluop  : std_logic_vector(2 downto 0);  	-- Alu operation
    alusel : std_logic_vector(1 downto 0);  	-- Alu result select
    aluadd : std_ulogic;
    alucin : std_ulogic;
    ldbp1, ldbp2 : std_ulogic;
    invop2 : std_ulogic;
    shcnt  : std_logic_vector(4 downto 0);  	-- shift count
    sari   : std_ulogic;				-- shift msb
    shleft : std_ulogic;				-- shift left/right
    ymsb   : std_ulogic;				-- shift left/right
    rd 	   : std_logic_vector(4 downto 0);
    jmpl   : std_ulogic;
    su     : std_ulogic;
    et     : std_ulogic;
    cwp    : cwptype;
    icc    : std_logic_vector(3 downto 0);
    mulstep: std_ulogic;            
    mul    : std_ulogic;            
    mac    : std_ulogic;
  end record;
  
  type memory_reg_type is record
    ctrl   : pipeline_ctrl_type;
    result : word;
    y      : word;
    icc    : std_logic_vector(3 downto 0);
    nalign : std_ulogic;
    dci	   : dc_in_type;
    werr   : std_ulogic;
    wcwp   : std_ulogic;
    irqen  : std_ulogic;
    irqen2 : std_ulogic;
    mac    : std_ulogic;
    divz   : std_ulogic;
    su     : std_ulogic;
    mul    : std_ulogic;
  end record;

  type exception_state is (run, trap, dsu1, dsu2);
  
  type exception_reg_type is record
    ctrl   : pipeline_ctrl_type;
    result : word;
    y      : word;
    icc    : std_logic_vector( 3 downto 0);
    annul_all : std_ulogic;
    data   : dcdtype;
    set    : std_logic_vector(0 downto 0);
    mexc   : std_ulogic;
    dci	   : dc_in_type;
    laddr  : std_logic_vector(1 downto 0);
    rstate : exception_state;
    npc    : std_logic_vector(2 downto 0);
    intack : std_ulogic;
    ipend  : std_ulogic;
    mac    : std_ulogic;
    debug  : std_ulogic;
    nerror : std_ulogic;
  end record;

  type dsu_registers is record
    tt      : std_logic_vector(7 downto 0);
    err     : std_ulogic;
    tbufcnt : std_logic_vector(7-1 downto 0);
    asi     : std_logic_vector(7 downto 0);
    crdy    : std_logic_vector(2 downto 1);  -- diag cache access ready
  end record;

  type irestart_register is record
    addr   : pctype;
    pwd    : std_ulogic;
  end record;
  
  type pwd_register_type is record
    pwd    : std_ulogic;
    error  : std_ulogic;
  end record;

  type special_register_type is record
    cwp    : cwptype;                             -- current window pointer
    icc    : std_logic_vector(3 downto 0);	  -- integer condition codes
    tt     : std_logic_vector(7 downto 0);	  -- trap type
    tba    : std_logic_vector(19 downto 0);	  -- trap base address
    wim    : std_logic_vector(8-1 downto 0);   -- window invalid mask
    pil    : std_logic_vector(3 downto 0);	  -- processor interrupt level
    ec     : std_ulogic;			   -- enable CP 
    ef     : std_ulogic;			   -- enable FP 
    ps     : std_ulogic;			   -- previous supervisor flag
    s      : std_ulogic;			   -- supervisor flag
    et     : std_ulogic;			   -- enable traps
    y      : word;
    asr18  : word;
    svt    : std_ulogic;			   -- enable traps
    dwt    : std_ulogic;			   -- disable write error trap
  end record;
  
  type write_reg_type is record
    s      : special_register_type;
    result : word;
    wa     : rfatype;
    wreg   : std_ulogic;
    except : std_ulogic;
  end record;

  type registers is record
    f  : fetch_reg_type;
    d  : decode_reg_type;
    a  : regacc_reg_type;
    e  : execute_reg_type;
    m  : memory_reg_type;
    x  : exception_reg_type;
    w  : write_reg_type;
  end record;

  type exception_type is record
    pri   : std_ulogic;
    ill   : std_ulogic;
    fpdis : std_ulogic;
    cpdis : std_ulogic;
    wovf  : std_ulogic;
    wunf  : std_ulogic;
    ticc  : std_ulogic;
  end record;

  type watchpoint_register is record
    addr    : std_logic_vector(31 downto 2);  -- watchpoint address
    mask    : std_logic_vector(31 downto 2);  -- watchpoint mask
    exec    : std_ulogic;			    -- trap on instruction
    load    : std_ulogic;			    -- trap on load
    store   : std_ulogic;			    -- trap on store
  end record;

  type watchpoint_registers is array (0 to 3) of watchpoint_register;

  constant wpr_none : watchpoint_register := (
	"000000000000000000000000000000", "000000000000000000000000000000", '0', '0', '0');

  function dbgexc(r  : registers; dbgi : l3_debug_in_type; trap : std_ulogic; tt : std_logic_vector(7 downto 0)) return std_ulogic is
    variable dmode : std_ulogic;
  begin
    dmode := '0';
    if (not r.x.ctrl.annul and trap) = '1' then
      if (((tt = "00" & TT_WATCH) and (dbgi.bwatch = '1')) or
          ((dbgi.bsoft = '1') and (tt = "10000001")) or
          (dbgi.btrapa = '1') or
          ((dbgi.btrape = '1') and not ((tt(5 downto 0) = TT_PRIV) or 
	    (tt(5 downto 0) = TT_FPDIS) or (tt(5 downto 0) = TT_WINOF) or
            (tt(5 downto 0) = TT_WINUF) or (tt(5 downto 4) = "01") or (tt(7) = '1'))) or 
          (((not r.w.s.et) and dbgi.berror) = '1')) then
        dmode := '1';
      end if;
    end if;
    return(dmode);
  end;
                    
  function dbgerr(r : registers; dbgi : l3_debug_in_type;
                  tt : std_logic_vector(7 downto 0))
  return std_ulogic is
    variable err : std_ulogic;
  begin
    err := not r.w.s.et;
    if (((dbgi.dbreak = '1') and (tt = ("00" & TT_WATCH))) or
        ((dbgi.bsoft = '1') and (tt = ("10000001")))) then
      err := '0';
    end if;
    return(err);
  end;
  
  procedure diagwr(r    : in registers;
                   dsur : in dsu_registers;
                   ir   : in irestart_register;
                   dbg  : in l3_debug_in_type;
                   wpr  : in watchpoint_registers;
                   s    : out special_register_type;
                   vwpr : out watchpoint_registers;
                   asi : out std_logic_vector(7 downto 0);
                   pc, npc  : out pctype;
                   tbufcnt : out std_logic_vector(7-1 downto 0);
                   wr : out std_ulogic;
                   addr : out std_logic_vector(9 downto 0);
                   data : out word;
                   fpcwr : out std_ulogic) is
  variable i : integer range 0 to 3;
  begin
    s := r.w.s; pc := r.f.pc; npc := ir.addr; wr := '0';
    vwpr := wpr; asi := dsur.asi; addr := "0000000000";
    data := dbg.ddata;
    tbufcnt := dsur.tbufcnt; fpcwr := '0';
      if (dbg.dsuen and dbg.denable and dbg.dwrite) = '1' then
        case dbg.daddr(23 downto 20) is
          when "0001" =>
            if (dbg.daddr(16) = '1') and true then -- trace buffer control reg
              tbufcnt := dbg.ddata(7-1 downto 0);
            end if;
          when "0011" => -- IU reg file
            if dbg.daddr(12) = '0' then
              wr := '1';
              addr := "0000000000";
              addr(8-1 downto 0) := dbg.daddr(8+1 downto 2);
            else  -- FPC
              fpcwr := '1';
            end if;
          when "0100" => -- IU special registers
            case dbg.daddr(7 downto 6) is
              when "00" => -- IU regs Y - TBUF ctrl reg
                case dbg.daddr(5 downto 2) is
                  when "0000" => -- Y
                    s.y := dbg.ddata;
                  when "0001" => -- PSR
                    s.cwp := dbg.ddata(3-1 downto 0);
                    s.icc := dbg.ddata(23 downto 20);
                    s.ec  := dbg.ddata(13);
                    if FPEN then s.ef := dbg.ddata(12); end if;
                    s.pil := dbg.ddata(11 downto 8);
                    s.s   := dbg.ddata(7);
                    s.ps  := dbg.ddata(6);
                    s.et  := dbg.ddata(5);
                  when "0010" => -- WIM
                    s.wim := dbg.ddata(8-1 downto 0);
                  when "0011" => -- TBR
                    s.tba := dbg.ddata(31 downto 12);
                    s.tt  := dbg.ddata(11 downto 4);
                  when "0100" => -- PC
                    pc := dbg.ddata(31 downto 2);
                  when "0101" => -- NPC
                    npc := dbg.ddata(31 downto 2);
                  when "0110" => --FSR
                    fpcwr := '1';
                  when "0111" => --CFSR
                  when "1001" => -- ASI reg
                    asi := dbg.ddata(7 downto 0);
                  --when "1001" => -- TBUF ctrl reg
                  --  tbufcnt := dbg.ddata(7-1 downto 0);
                  when others =>
                end case;
              when "01" => -- ASR16 - ASR31
		case dbg.daddr(5 downto 2) is
		when "0001" =>	-- %ASR17
	    	  s.dwt := dbg.ddata(14);
	    	  s.svt := dbg.ddata(13);
		when "0010" =>	-- %ASR18
		  if false then s.asr18 := dbg.ddata; end if;
		when "1000" => 		-- %ASR24 - %ASR31
                  vwpr(0).addr := dbg.ddata(31 downto 2);
                  vwpr(0).exec := dbg.ddata(0); 
		when "1001" =>
                  vwpr(0).mask := dbg.ddata(31 downto 2);
                  vwpr(0).load := dbg.ddata(1);
                  vwpr(0).store := dbg.ddata(0);              
		when "1010" =>
                  vwpr(1).addr := dbg.ddata(31 downto 2);
                  vwpr(1).exec := dbg.ddata(0); 
		when "1011" =>
                  vwpr(1).mask := dbg.ddata(31 downto 2);
                  vwpr(1).load := dbg.ddata(1);
                  vwpr(1).store := dbg.ddata(0);              
		when "1100" =>
                  vwpr(2).addr := dbg.ddata(31 downto 2);
                  vwpr(2).exec := dbg.ddata(0); 
		when "1101" =>
                  vwpr(2).mask := dbg.ddata(31 downto 2);
                  vwpr(2).load := dbg.ddata(1);
                  vwpr(2).store := dbg.ddata(0);              
		when "1110" =>
                  vwpr(3).addr := dbg.ddata(31 downto 2);
                  vwpr(3).exec := dbg.ddata(0); 
		when "1111" => -- 
                  vwpr(3).mask := dbg.ddata(31 downto 2);
                  vwpr(3).load := dbg.ddata(1);
                  vwpr(3).store := dbg.ddata(0);              
		when others => -- 
		end case;
-- disabled due to bug in XST
--                  i := conv_integer(dbg.daddr(4 downto 3)); 
--                  if dbg.daddr(2) = '0' then
--                    vwpr(i).addr := dbg.ddata(31 downto 2);
--                    vwpr(i).exec := dbg.ddata(0); 
--                  else
--                    vwpr(i).mask := dbg.ddata(31 downto 2);
--                    vwpr(i).load := dbg.ddata(1);
--                    vwpr(i).store := dbg.ddata(0);              
--                  end if;                    
              when others =>
            end case;
          when others =>
        end case;
      end if;
  end;

  function asr17_gen ( r : in registers) return word is
  variable asr17 : word;
  variable fpu2 : integer range 0 to 3;
  begin
    asr17 := "00000000000000000000000000000000";    
    asr17(31 downto 28) := conv_std_logic_vector(index, 4);
    if (clk2x > 8) then
      asr17(16 downto 15) := conv_std_logic_vector(clk2x-8, 2);
      asr17(17) := '1'; 
    elsif (clk2x > 0) then
      asr17(16 downto 15) := conv_std_logic_vector(clk2x, 2);
    end if;
    asr17(14) := r.w.s.dwt;
    if svt = 1 then asr17(13) := r.w.s.svt; end if;
    if lddel = 2 then asr17(12) := '1'; end if;
    if (fpu > 0) and (fpu < 8) then fpu2 := 1;
    elsif (fpu >= 8) and (fpu < 15) then fpu2 := 3;                          
    elsif fpu = 15 then fpu2 := 2;
    else fpu2 := 0; end if; 
    asr17(11 downto 10) := conv_std_logic_vector(fpu2, 2);                       
    if mac = 1 then asr17(9) := '1'; end if;
    if 2 /= 0 then asr17(8) := '1'; end if;
    asr17(7 downto 5) := conv_std_logic_vector(nwp, 3);                       
    asr17(4 downto 0) := conv_std_logic_vector(8-1, 5);       
    return(asr17);
  end;

  procedure diagread(dbgi   : in l3_debug_in_type;
                     r      : in registers;
                     dsur   : in dsu_registers;
                     ir     : in irestart_register;
                     wpr    : in watchpoint_registers;
                     dco   : in  dcache_out_type;                          
                     tbufo  : in tracebuf_out_type;
                     data : out word) is
    variable cwp : std_logic_vector(4 downto 0);
    variable rd : std_logic_vector(4 downto 0);
    variable i : integer range 0 to 3;    
  begin
    data := "00000000000000000000000000000000"; cwp := "00000";
    cwp(3-1 downto 0) := r.w.s.cwp;
      case dbgi.daddr(22 downto 20) is
        when "001" => -- trace buffer
	  if true then
            if dbgi.daddr(16) = '1' then -- trace buffer control reg
              if true then data(7-1 downto 0) := dsur.tbufcnt; end if;
            else
              case dbgi.daddr(3 downto 2) is
              when "00" => data := tbufo.data(127 downto 96);
              when "01" => data := tbufo.data(95 downto 64);
              when "10" => data := tbufo.data(63 downto 32);
              when others => data := tbufo.data(31 downto 0);
              end case;
            end if;
          end if;
        when "011" => -- IU reg file
          if dbgi.daddr(12) = '0' then
            data := rfo.data1(31 downto 0); 
            if (dbgi.daddr(11) = '1') and (is_fpga(fabtech) = 0) then 
	      data := rfo.data2(31 downto 0);
	    end if;
          else data := fpo.dbg.data; end if;
        when "100" => -- IU regs
          case dbgi.daddr(7 downto 6) is
            when "00" => -- IU regs Y - TBUF ctrl reg
              case dbgi.daddr(5 downto 2) is
                when "0000" =>
                  data := r.w.s.y;
                when "0001" =>
                  data := conv_std_logic_vector(15, 4) & conv_std_logic_vector(3, 4) &
                          r.w.s.icc & "000000" & r.w.s.ec & r.w.s.ef & r.w.s.pil &
                          r.w.s.s & r.w.s.ps & r.w.s.et & cwp;
                when "0010" =>
                  data(8-1 downto 0) := r.w.s.wim;
                when "0011" =>
                  data := r.w.s.tba & r.w.s.tt & "0000";
                when "0100" =>
                  data(31 downto 2) := r.f.pc;
                when "0101" =>
                  data(31 downto 2) := ir.addr;
                when "0110" => -- FSR
                  data := fpo.dbg.data;
                when "0111" => -- CPSR
                when "1000" => -- TT reg
                  data(12 downto 4) := dsur.err & dsur.tt;
                when "1001" => -- ASI reg
                  data(7 downto 0) := dsur.asi;
                when others =>
              end case;
            when "01" =>
              if dbgi.daddr(5) = '0' then -- %ASR17
                if dbgi.daddr(4 downto 2) = "001" then -- %ASR17
		  data := asr17_gen(r);
		elsif false and  dbgi.daddr(4 downto 2) = "010" then -- %ASR18
		  data := r.w.s.asr18;
		end if;
              else  -- %ASR24 - %ASR31
                i := conv_integer(dbgi.daddr(4 downto 3));                                           -- 
                if dbgi.daddr(2) = '0' then
                  data(31 downto 2) := wpr(i).addr;
                  data(0) := wpr(i).exec;
                else
                  data(31 downto 2) := wpr(i).mask;
                  data(1) := wpr(i).load;
                  data(0) := wpr(i).store; 
                end if;
              end if;
            when others =>
          end case;
        when "111" =>
          data := r.x.data(conv_integer(r.x.set));
        when others =>
      end case;
  end;
  

  procedure itrace(r    : in registers;
                   dsur : in dsu_registers;
                   vdsu : in dsu_registers;
                   res  : in word;
                   exc  : in std_ulogic;
                   dbgi : in l3_debug_in_type;
                   error : in std_ulogic;
                   trap  : in std_ulogic;                          
                   tbufcnt : out std_logic_vector(7-1 downto 0); 
                   di  : out tracebuf_in_type) is
  variable meminst : std_ulogic;
  begin
    di.addr := (others => '0'); di.data := (others => '0');
    di.enable := '0'; di.write := (others => '0');
    tbufcnt := vdsu.tbufcnt;
    meminst := r.x.ctrl.inst(31) and r.x.ctrl.inst(30);
    if true then
      di.addr(7-1 downto 0) := dsur.tbufcnt;
      di.data(127) := '0';
      di.data(126) := not r.x.ctrl.pv;
      di.data(125 downto 96) := dbgi.timer(29 downto 0);
      di.data(95 downto 64) := res;
      di.data(63 downto 34) := r.x.ctrl.pc(31 downto 2);
      di.data(33) := trap;
      di.data(32) := error;
      di.data(31 downto 0) := r.x.ctrl.inst;
      if (dbgi.tenable = '0') or (r.x.rstate = dsu2) then
        if ((dbgi.dsuen and dbgi.denable) = '1') and (dbgi.daddr(23 downto 20) & dbgi.daddr(16) = "00010") then
          di.enable := '1'; 
          di.addr(7-1 downto 0) := dbgi.daddr(7-1+4 downto 4);
          if dbgi.dwrite = '1' then            
            case dbgi.daddr(3 downto 2) is
              when "00" => di.write(3) := '1';
              when "01" => di.write(2) := '1';
              when "10" => di.write(1) := '1';
              when others => di.write(0) := '1';
            end case;
            di.data := dbgi.ddata & dbgi.ddata & dbgi.ddata & dbgi.ddata;
          end if;
        end if;
      elsif (not r.x.ctrl.annul and (r.x.ctrl.pv or meminst) and not r.x.debug) = '1' then        
        di.enable := '1'; di.write := (others => '1');
        tbufcnt := dsur.tbufcnt + 1;
      end if;
      di.diag := dco.testen & "000";
      if dco.scanen = '1' then di.enable := '0'; end if;
    end if;
  end;

  procedure dbg_cache(holdn    : in std_ulogic;
                      dbgi     :  in l3_debug_in_type;
                      r        : in registers;
                      dsur     : in dsu_registers;
                      mresult  : in word;
                      dci      : in dc_in_type;
                      mresult2 : out word;
                      dci2     : out dc_in_type
                      ) is
  begin
    mresult2 := mresult; dci2 := dci; dci2.dsuen := '0'; 
    if true then
      if r.x.rstate = dsu2 then
        dci2.asi := dsur.asi;
        if (dbgi.daddr(22 downto 20) = "111") and (dbgi.dsuen = '1') then
          dci2.dsuen := (dbgi.denable or r.m.dci.dsuen) and not dsur.crdy(2);
          dci2.enaddr := dbgi.denable;
          dci2.size := "10"; dci2.read := '1'; dci2.write := '0';
          if (dbgi.denable and not r.m.dci.enaddr) = '1' then            
            mresult2 := (others => '0'); mresult2(19 downto 2) := dbgi.daddr(19 downto 2);
          else
            mresult2 := dbgi.ddata;            
          end if;
          if dbgi.dwrite = '1' then
            dci2.read := '0'; dci2.write := '1';
          end if;
        end if;
      end if;
    end if;
  end;
    
  procedure fpexack(r : in registers; fpexc : out std_ulogic) is
  begin
    fpexc := '0';
    if FPEN then 
      if r.x.ctrl.tt = TT_FPEXC then fpexc := '1'; end if;
    end if;
  end;

  procedure diagrdy(denable : in std_ulogic;
                    dsur : in dsu_registers;
                    dci   : in dc_in_type;
                    mds : in std_ulogic;
                    ico : in icache_out_type;
                    crdy : out std_logic_vector(2 downto 1)) is                   
  begin
    crdy := dsur.crdy(1) & '0';    
    if dci.dsuen = '1' then
      case dsur.asi(4 downto 0) is
        when ASI_ITAG | ASI_IDATA | ASI_UINST | ASI_SINST =>
          crdy(2) := ico.diagrdy and not dsur.crdy(2);
        when ASI_DTAG | ASI_MMUSNOOP_DTAG | ASI_DDATA | ASI_UDATA | ASI_SDATA =>
          crdy(1) := not denable and dci.enaddr and not dsur.crdy(1);
        when others =>
          crdy(2) := dci.enaddr and denable;
      end case;
    end if;
  end;

  
  signal r, rin : registers;
  signal wpr, wprin : watchpoint_registers;
  signal dsur, dsuin : dsu_registers;
  signal ir, irin : irestart_register;
  signal rp, rpin : pwd_register_type;

-- execute stage operations

  constant EXE_AND   : std_logic_vector(2 downto 0) := "000";
  constant EXE_XOR   : std_logic_vector(2 downto 0) := "001"; -- must be equal to EXE_PASS2
  constant EXE_OR    : std_logic_vector(2 downto 0) := "010";
  constant EXE_XNOR  : std_logic_vector(2 downto 0) := "011";
  constant EXE_ANDN  : std_logic_vector(2 downto 0) := "100";
  constant EXE_ORN   : std_logic_vector(2 downto 0) := "101";
  constant EXE_DIV   : std_logic_vector(2 downto 0) := "110";

  constant EXE_PASS1 : std_logic_vector(2 downto 0) := "000";
  constant EXE_PASS2 : std_logic_vector(2 downto 0) := "001";
  constant EXE_STB   : std_logic_vector(2 downto 0) := "010";
  constant EXE_STH   : std_logic_vector(2 downto 0) := "011";
  constant EXE_ONES  : std_logic_vector(2 downto 0) := "100";
  constant EXE_RDY   : std_logic_vector(2 downto 0) := "101";
  constant EXE_SPR   : std_logic_vector(2 downto 0) := "110";
  constant EXE_LINK  : std_logic_vector(2 downto 0) := "111";

  constant EXE_SLL   : std_logic_vector(2 downto 0) := "001";
  constant EXE_SRL   : std_logic_vector(2 downto 0) := "010";
  constant EXE_SRA   : std_logic_vector(2 downto 0) := "100";

  constant EXE_NOP   : std_logic_vector(2 downto 0) := "000";

-- EXE result select

  constant EXE_RES_ADD   : std_logic_vector(1 downto 0) := "00";
  constant EXE_RES_SHIFT : std_logic_vector(1 downto 0) := "01";
  constant EXE_RES_LOGIC : std_logic_vector(1 downto 0) := "10";
  constant EXE_RES_MISC  : std_logic_vector(1 downto 0) := "11";

-- Load types

  constant SZBYTE    : std_logic_vector(1 downto 0) := "00";
  constant SZHALF    : std_logic_vector(1 downto 0) := "01";
  constant SZWORD    : std_logic_vector(1 downto 0) := "10";
  constant SZDBL     : std_logic_vector(1 downto 0) := "11";

-- calculate register file address

  procedure regaddr(cwp : std_logic_vector; reg : std_logic_vector(4 downto 0);
	 rao : out rfatype) is
  variable ra : rfatype;
  constant globals : std_logic_vector(8-5  downto 0) := 
	conv_std_logic_vector(8, 8-4);
  begin
    ra := (others => '0'); ra(4 downto 0) := reg;
    if reg(4 downto 3) = "00" then ra(8 -1 downto 4) := globals;
    else
      ra(3+3 downto 4) := cwp + ra(4);
      if ra(8-1 downto 4) = globals then
        ra(8-1 downto 4) := (others => '0');
      end if;
    end if;
    rao := ra;
  end;

-- branch adder

  function branch_address(inst : word; pc : pctype) return std_logic_vector is
  variable baddr, caddr, tmp : pctype;
  begin
    caddr := (others => '0'); caddr(31 downto 2) := inst(29 downto 0);
    caddr(31 downto 2) := caddr(31 downto 2) + pc(31 downto 2);
    baddr := (others => '0'); baddr(31 downto 24) := (others => inst(21)); 
    baddr(23 downto 2) := inst(21 downto 0);
    baddr(31 downto 2) := baddr(31 downto 2) + pc(31 downto 2);
    if inst(30) = '1' then tmp := caddr; else tmp := baddr; end if;
    return(tmp);
  end;

-- evaluate branch condition

  function branch_true(icc : std_logic_vector(3 downto 0); inst : word) 
	return std_ulogic is
  variable n, z, v, c, branch : std_ulogic;
  begin
    n := icc(3); z := icc(2); v := icc(1); c := icc(0);
    case inst(27 downto 25) is
    when "000" =>  branch := inst(28) xor '0';			-- bn, ba
    when "001" =>  branch := inst(28) xor z;      		-- be, bne
    when "010" =>  branch := inst(28) xor (z or (n xor v));     -- ble, bg
    when "011" =>  branch := inst(28) xor (n xor v); 	        -- bl, bge
    when "100" =>  branch := inst(28) xor (c or z);   	        -- bleu, bgu
    when "101" =>  branch := inst(28) xor c;		        -- bcs, bcc 
    when "110" =>  branch := inst(28) xor n;		        -- bneg, bpos
    when others => branch := inst(28) xor v;		        -- bvs, bvc   
    end case;
    return(branch);
  end;

-- detect RETT instruction in the pipeline and set the local psr.su and psr.et

  procedure su_et_select(r : in registers; xc_ps, xc_s, xc_et : in std_ulogic;
		       su, et : out std_ulogic) is
  begin
   if ((r.a.ctrl.rett or r.e.ctrl.rett or r.m.ctrl.rett or r.x.ctrl.rett) = '1')
     and (r.x.annul_all = '0')
   then su := xc_ps; et := '1';
   else su := xc_s; et := xc_et; end if;
  end;

-- detect watchpoint trap

  function wphit(r : registers; wpr : watchpoint_registers; debug : l3_debug_in_type)
    return std_ulogic is
  variable exc : std_ulogic;
  begin
    exc := '0';
    for i in 1 to NWP loop
      if ((wpr(i-1).exec and r.a.ctrl.pv and not r.a.ctrl.annul) = '1') then
         if (((wpr(i-1).addr xor r.a.ctrl.pc(31 downto 2)) and wpr(i-1).mask) = "000000000000000000000000000000") then
           exc := '1';
	 end if;
      end if;
    end loop;

   if true then
     if (debug.dsuen and not r.a.ctrl.annul) = '1' then
       exc := exc or (r.a.ctrl.pv and ((debug.dbreak and debug.bwatch) or r.a.step));
     end if;
   end if;
    return(exc);
  end;

-- 32-bit shifter

  function shift3(r : registers; aluin1, aluin2 : word) return word is
  variable shiftin : unsigned(63 downto 0);
  variable shiftout : unsigned(63 downto 0);
  variable cnt : natural range 0 to 31;
  begin

    cnt := conv_integer(r.e.shcnt);
    if r.e.shleft = '1' then
      shiftin(30 downto 0) := (others => '0');
      shiftin(63 downto 31) := '0' & unsigned(aluin1);
    else
      shiftin(63 downto 32) := (others => r.e.sari);
      shiftin(31 downto 0) := unsigned(aluin1);
    end if;
    shiftout := SHIFT_RIGHT(shiftin, cnt);
    return(std_logic_vector(shiftout(31 downto 0)));
     
  end;

  function shift2(r : registers; aluin1, aluin2 : word) return word is
  variable ushiftin : unsigned(31 downto 0);
  variable sshiftin : signed(32 downto 0);
  variable cnt : natural range 0 to 31;
  variable resleft, resright : word;
  begin

    cnt := conv_integer(r.e.shcnt);
    ushiftin := unsigned(aluin1);
    sshiftin := signed('0' & aluin1);
    if r.e.shleft = '1' then
      resleft := std_logic_vector(SHIFT_LEFT(ushiftin, cnt));
      return(resleft);
    else
      if r.e.sari = '1' then sshiftin(32) := aluin1(31); end if;
      sshiftin := SHIFT_RIGHT(sshiftin, cnt);
      resright := std_logic_vector(sshiftin(31 downto 0));
      return(resright);
--      else 
--	ushiftin := SHIFT_RIGHT(ushiftin, cnt);
--        return(std_logic_vector(ushiftin));
--      end if;
    end if;
     
  end;

  function shift(r : registers; aluin1, aluin2 : word;
	         shiftcnt : std_logic_vector(4 downto 0); sari : std_ulogic ) return word is
  variable shiftin : std_logic_vector(63 downto 0);
  begin
    shiftin := "00000000000000000000000000000000" & aluin1;
    if r.e.shleft = '1' then
      shiftin(31 downto 0) := "00000000000000000000000000000000"; shiftin(63 downto 31) := '0' & aluin1;
    else shiftin(63 downto 32) := (others => sari); end if;
    if shiftcnt (4) = '1' then shiftin(47 downto 0) := shiftin(63 downto 16); end if;
    if shiftcnt (3) = '1' then shiftin(39 downto 0) := shiftin(47 downto 8); end if;
    if shiftcnt (2) = '1' then shiftin(35 downto 0) := shiftin(39 downto 4); end if;
    if shiftcnt (1) = '1' then shiftin(33 downto 0) := shiftin(35 downto 2); end if;
    if shiftcnt (0) = '1' then shiftin(31 downto 0) := shiftin(32 downto 1); end if;
    return(shiftin(31 downto 0));
  end;

-- Check for illegal and privileged instructions

procedure exception_detect(r : registers; wpr : watchpoint_registers; dbgi : l3_debug_in_type;
        trapin : in std_ulogic; ttin : in std_logic_vector(5 downto 0); 
	trap : out std_ulogic; tt : out std_logic_vector(5 downto 0)) is
variable illegal_inst, privileged_inst : std_ulogic;
variable cp_disabled, fp_disabled, fpop : std_ulogic;
variable op : std_logic_vector(1 downto 0);
variable op2 : std_logic_vector(2 downto 0);
variable op3 : std_logic_vector(5 downto 0);
variable rd  : std_logic_vector(4 downto 0);
variable inst : word;
variable wph : std_ulogic;
begin
  inst := r.a.ctrl.inst; trap := trapin; tt := ttin;
  if r.a.ctrl.annul = '0' then
    op  := inst(31 downto 30); op2 := inst(24 downto 22);
    op3 := inst(24 downto 19); rd  := inst(29 downto 25);
    illegal_inst := '0'; privileged_inst := '0'; cp_disabled := '0'; 
    fp_disabled := '0'; fpop := '0';
    case op is
    when CALL => null;
    when FMT2 =>
      case op2 is
      when SETHI | BICC => null;
      when FBFCC => 
	if FPEN then fp_disabled := not r.w.s.ef; else fp_disabled := '1'; end if;
      when CBCCC =>
	if (not false) or (r.w.s.ec = '0') then cp_disabled := '1'; end if;
      when others => illegal_inst := '1';
      end case;
    when FMT3 =>
      case op3 is
      when IAND | ANDCC | ANDN | ANDNCC | IOR | ORCC | ORN | ORNCC | IXOR |
        XORCC | IXNOR | XNORCC | ISLL | ISRL | ISRA | MULSCC | IADD | ADDX |
	ADDCC | ADDXCC | ISUB | SUBX | SUBCC | SUBXCC | FLUSH | JMPL | TICC | 
	SAVE | RESTORE | RDY => null;
      when TADDCC | TADDCCTV | TSUBCC | TSUBCCTV => 
	if notag = 1 then illegal_inst := '1'; end if;
      when UMAC | SMAC => 
	if not false then illegal_inst := '1'; end if;
      when UMUL | SMUL | UMULCC | SMULCC => 
	if not true then illegal_inst := '1'; end if;
      when UDIV | SDIV | UDIVCC | SDIVCC => 
	if not true then illegal_inst := '1'; end if;
      when RETT => illegal_inst := r.a.et; privileged_inst := not r.a.su;
      when RDPSR | RDTBR | RDWIM => privileged_inst := not r.a.su;
      when WRY  => null;
      when WRPSR => 
	privileged_inst := not r.a.su; 
      when WRWIM | WRTBR  => privileged_inst := not r.a.su;
      when FPOP1 | FPOP2 => 
	if FPEN then fp_disabled := not r.w.s.ef; fpop := '1';
	else fp_disabled := '1'; fpop := '0'; end if;
      when CPOP1 | CPOP2 =>
	if (not false) or (r.w.s.ec = '0') then cp_disabled := '1'; end if;
      when others => illegal_inst := '1';
      end case;
    when others =>	-- LDST
      case op3 is
      when LDD | ISTD => illegal_inst := rd(0);	-- trap if odd destination register
      when LD | LDUB | LDSTUB | LDUH | LDSB | LDSH | ST | STB | STH | SWAP =>
	null;
      when LDDA | STDA =>
	illegal_inst := inst(13) or rd(0); privileged_inst := not r.a.su;
      when LDA | LDUBA| LDSTUBA | LDUHA | LDSBA | LDSHA | STA | STBA | STHA |
	   SWAPA => 
	illegal_inst := inst(13); privileged_inst := not r.a.su;
      when LDDF | STDF | LDF | LDFSR | STF | STFSR => 
	if FPEN then fp_disabled := not r.w.s.ef;
	else fp_disabled := '1'; end if;
      when STDFQ => 
	privileged_inst := not r.a.su; 
	if (not FPEN) or (r.w.s.ef = '0') then fp_disabled := '1'; end if;
      when STDCQ => 
	privileged_inst := not r.a.su;
	if (not false) or (r.w.s.ec = '0') then cp_disabled := '1'; end if;
      when LDC | LDCSR | LDDC | STC | STCSR | STDC => 
	if (not false) or (r.w.s.ec = '0') then cp_disabled := '1'; end if;
      when others => illegal_inst := '1';
      end case;
    end case;

    wph := wphit(r, wpr, dbgi);
    
    trap := '1';
    if r.a.ctrl.trap = '1' then tt := TT_IAEX;
    elsif privileged_inst = '1' then tt := TT_PRIV; 
    elsif illegal_inst = '1' then tt := TT_IINST;
    elsif fp_disabled = '1' then tt := TT_FPDIS;
    elsif cp_disabled = '1' then tt := TT_CPDIS;
    elsif wph = '1' then tt := TT_WATCH;
    elsif r.a.wovf= '1' then tt := TT_WINOF;
    elsif r.a.wunf= '1' then tt := TT_WINUF;
    elsif r.a.ticc= '1' then tt := TT_TICC;
    else trap := '0'; tt:= (others => '0'); end if;
  end if;
end;

-- instructions that write the condition codes (psr.icc)

procedure wicc_y_gen(inst : word; wicc, wy : out std_ulogic) is
begin
  wicc := '0'; wy := '0';
  if inst(31 downto 30) = FMT3 then
    case inst(24 downto 19) is
    when SUBCC | TSUBCC | TSUBCCTV | ADDCC | ANDCC | ORCC | XORCC | ANDNCC |
	 ORNCC | XNORCC | TADDCC | TADDCCTV | ADDXCC | SUBXCC | WRPSR => 
      wicc := '1';
    when WRY =>
      if r.d.inst(conv_integer(r.d.set))(29 downto 25) = "00000" then wy := '1'; end if;
    when MULSCC =>
      wicc := '1'; wy := '1';
    when  UMAC | SMAC  =>
      if false then wy := '1'; end if;
    when UMULCC | SMULCC => 
      if true and (((mulo.nready = '1') and (r.d.cnt /= "00")) or (0 /= 0)) then
        wicc := '1'; wy := '1';
      end if;
    when UMUL | SMUL => 
      if true and (((mulo.nready = '1') and (r.d.cnt /= "00")) or (0 /= 0)) then
        wy := '1';
      end if;
    when UDIVCC | SDIVCC => 
      if true and (divo.nready = '1') and (r.d.cnt /= "00") then
        wicc := '1';
      end if;
    when others =>
    end case;
  end if;
end;

-- select cwp 

procedure cwp_gen(r, v : registers; annul, wcwp : std_ulogic; ncwp : cwptype;
		  cwp : out cwptype) is
begin
  if (r.x.rstate = trap) or (r.x.rstate = dsu2) or (rstn = '0') then cwp := v.w.s.cwp;
  elsif (wcwp = '1') and (annul = '0') then cwp := ncwp;
  elsif r.m.wcwp = '1' then cwp := r.m.result(3-1 downto 0);
  else cwp := r.d.cwp; end if;
end;

-- generate wcwp in ex stage

procedure cwp_ex(r : in  registers; wcwp : out std_ulogic) is
begin
  if (r.e.ctrl.inst(31 downto 30) = FMT3) and 
     (r.e.ctrl.inst(24 downto 19) = WRPSR)
  then wcwp := not r.e.ctrl.annul; else wcwp := '0'; end if;
end;

-- generate next cwp & window under- and overflow traps

procedure cwp_ctrl(r : in registers; xc_wim : in std_logic_vector(8-1 downto 0);
	inst : word; de_cwp : out cwptype; wovf_exc, wunf_exc, wcwp : out std_ulogic) is
variable op : std_logic_vector(1 downto 0);
variable op3 : std_logic_vector(5 downto 0);
variable wim : word;
variable ncwp : cwptype;
begin
  op := inst(31 downto 30); op3 := inst(24 downto 19); 
  wovf_exc := '0'; wunf_exc := '0'; wim := (others => '0'); 
  wim(8-1 downto 0) := xc_wim; ncwp := r.d.cwp; wcwp := '0';

  if (op = FMT3) and ((op3 = RETT) or (op3 = RESTORE) or (op3 = SAVE)) then
    wcwp := '1';
    if (op3 = SAVE) then
      if (not true) and (r.d.cwp = "000") then ncwp := "111";
      else ncwp := r.d.cwp - 1 ; end if;
    else
      if (not true) and (r.d.cwp = "111") then ncwp := "000";
      else ncwp := r.d.cwp + 1; end if;
    end if;
    if wim(conv_integer(ncwp)) = '1' then
      if op3 = SAVE then wovf_exc := '1'; else wunf_exc := '1'; end if;
    end if;
  end if;
  de_cwp := ncwp;
end;

-- generate register read address 1

procedure rs1_gen(r : registers; inst : word;  rs1 : out std_logic_vector(4 downto 0);
	rs1mod : out std_ulogic) is
variable op : std_logic_vector(1 downto 0);
variable op3 : std_logic_vector(5 downto 0);
begin
  op := inst(31 downto 30); op3 := inst(24 downto 19); 
  rs1 := inst(18 downto 14); rs1mod := '0';
  if (op = LDST) then
    if ((r.d.cnt = "01") and ((op3(2) and not op3(3)) = '1')) or
        (r.d.cnt = "10") 
    then rs1mod := '1'; rs1 := inst(29 downto 25); end if;
    if ((r.d.cnt = "10") and (op3(3 downto 0) = "0111")) then
      rs1(0) := '1';
    end if;
  end if;
end;

-- load/icc interlock detection

  procedure lock_gen(r : registers; rs2, rd : std_logic_vector(4 downto 0);
	rfa1, rfa2, rfrd : rfatype; inst : word; fpc_lock, mulinsn, divinsn : std_ulogic;
        lldcheck1, lldcheck2, lldlock, lldchkra, lldchkex : out std_ulogic) is
  variable op : std_logic_vector(1 downto 0);
  variable op2 : std_logic_vector(2 downto 0);
  variable op3 : std_logic_vector(5 downto 0);
  variable cond : std_logic_vector(3 downto 0);
  variable rs1  : std_logic_vector(4 downto 0);
  variable i, ldcheck1, ldcheck2, ldchkra, ldchkex, ldcheck3 : std_ulogic;
  variable ldlock, icc_check, bicc_hold, chkmul, y_check : std_ulogic;
  variable lddlock : boolean;
  begin
    op := inst(31 downto 30); op3 := inst(24 downto 19); 
    op2 := inst(24 downto 22); cond := inst(28 downto 25); 
    rs1 := inst(18 downto 14); lddlock := false; i := inst(13);
    ldcheck1 := '0'; ldcheck2 := '0'; ldcheck3 := '0'; ldlock := '0';
    ldchkra := '1'; ldchkex := '1'; icc_check := '0'; bicc_hold := '0';
    y_check := '0';

    if (r.d.annul = '0') then
      case op is
      when FMT2 =>
	if (op2 = BICC) and (cond(2 downto 0) /= "000") then 
	  icc_check := '1';
	end if;
      when FMT3 =>
        ldcheck1 := '1'; ldcheck2 := not i;
        case op3 is
	when TICC =>
	  if (cond(2 downto 0) /= "000") then icc_check := '1'; end if;
        when RDY => 
          ldcheck1 := '0'; ldcheck2 := '0';
	  if false then y_check := '1'; end if;
        when RDWIM | RDTBR => 
          ldcheck1 := '0'; ldcheck2 := '0';
        when RDPSR => 
          ldcheck1 := '0'; ldcheck2 := '0'; icc_check := '1';
	  if true then icc_check := '1'; end if;
--	when ADDX | ADDXCC | SUBX | SUBXCC =>
--	  if true then icc_check := '1'; end if;
	when SDIV | SDIVCC | UDIV | UDIVCC =>
	  if true then y_check := '1'; end if;
        when FPOP1 | FPOP2 => ldcheck1:= '0'; ldcheck2 := '0';
        when others => 
        end case;
      when LDST =>
        ldcheck1 := '1'; ldchkra := '0';
	case r.d.cnt is
	when "00" =>
          if (lddel = 2) and (op3(2) = '1') then ldcheck3 := '1'; end if; 
          ldcheck2 := not i; ldchkra := '1';
	when "01" => ldcheck2 := not i;
	when others => ldchkex := '0';
        end case;
        if  (op3(2 downto 0) = "011") then lddlock := true; end if;
      when others => null;
      end case;
    end if;

    if true or true then 
      chkmul := mulinsn;
      bicc_hold := bicc_hold or (icc_check and r.m.ctrl.wicc and (r.m.ctrl.cnt(0) or r.m.mul));
    else chkmul := '0'; end if;
    if true then 
      bicc_hold := bicc_hold or (y_check and (r.a.ctrl.wy or r.e.ctrl.wy));
      chkmul := chkmul or divinsn;
    end if;

    bicc_hold := bicc_hold or (icc_check and (r.a.ctrl.wicc or r.e.ctrl.wicc));

    if (((r.a.ctrl.ld or chkmul) and r.a.ctrl.wreg and ldchkra) = '1') and
       (((ldcheck1 = '1') and (r.a.ctrl.rd = rfa1)) or
        ((ldcheck2 = '1') and (r.a.ctrl.rd = rfa2)) or
        ((ldcheck3 = '1') and (r.a.ctrl.rd = rfrd)))
    then ldlock := '1'; end if;

    if (((r.e.ctrl.ld or r.e.mac) and r.e.ctrl.wreg and ldchkex) = '1') and 
        ((lddel = 2) or (false and (r.e.mac = '1')) or ((0 = 3) and (r.e.mul = '1'))) and
       (((ldcheck1 = '1') and (r.e.ctrl.rd = rfa1)) or
        ((ldcheck2 = '1') and (r.e.ctrl.rd = rfa2)))
    then ldlock := '1'; end if;

    ldlock := ldlock or bicc_hold or fpc_lock;

    lldcheck1 := ldcheck1; lldcheck2:= ldcheck2; lldlock := ldlock;
    lldchkra := ldchkra; lldchkex := ldchkex;
  end;

  procedure fpbranch(inst : in word; fcc  : in std_logic_vector(1 downto 0);
                      branch : out std_ulogic) is
  variable cond : std_logic_vector(3 downto 0);
  variable fbres : std_ulogic;
  begin
    cond := inst(28 downto 25);
    case cond(2 downto 0) is
      when "000" => fbres := '0';			-- fba, fbn
      when "001" => fbres := fcc(1) or fcc(0);
      when "010" => fbres := fcc(1) xor fcc(0);
      when "011" => fbres := fcc(0);
      when "100" => fbres := (not fcc(1)) and fcc(0);
      when "101" => fbres := fcc(1);
      when "110" => fbres := fcc(1) and not fcc(0);
      when others => fbres := fcc(1) and fcc(0);
    end case;
    branch := cond(3) xor fbres;     
  end;

-- PC generation

  procedure ic_ctrl(r : registers; inst : word; annul_all, ldlock, branch_true, 
	fbranch_true, cbranch_true, fccv, cccv : in std_ulogic; 
	cnt : out std_logic_vector(1 downto 0); 
	de_pc : out pctype; de_branch, ctrl_annul, de_annul, jmpl_inst, inull, 
	de_pv, ctrl_pv, de_hold_pc, ticc_exception, rett_inst, mulstart,
	divstart : out std_ulogic) is
  variable op : std_logic_vector(1 downto 0);
  variable op2 : std_logic_vector(2 downto 0);
  variable op3 : std_logic_vector(5 downto 0);
  variable cond : std_logic_vector(3 downto 0);
  variable hold_pc, annul_current, annul_next, branch, annul, pv : std_ulogic;
  variable de_jmpl : std_ulogic;
  begin
    branch := '0'; annul_next := '0'; annul_current := '0'; pv := '1';
    hold_pc := '0'; ticc_exception := '0'; rett_inst := '0';
    op := inst(31 downto 30); op3 := inst(24 downto 19); 
    op2 := inst(24 downto 22); cond := inst(28 downto 25); 
    annul := inst(29); de_jmpl := '0'; cnt := "00";
    mulstart := '0'; divstart := '0'; 
    if r.d.annul = '0' then
      case inst(31 downto 30) is
      when CALL =>
        branch := '1';
	if r.d.inull = '1' then 
	  hold_pc := '1'; annul_current := '1';
 	end if;
      when FMT2 =>
        if (op2 = BICC) or (FPEN and (op2 = FBFCC)) or (false and (op2 = CBCCC)) then
          if (FPEN and (op2 = FBFCC)) then 
	    branch := fbranch_true;
	    if fccv /= '1' then hold_pc := '1'; annul_current := '1'; end if;
          elsif (false and (op2 = CBCCC)) then 
	    branch := cbranch_true;
	    if cccv /= '1' then hold_pc := '1'; annul_current := '1'; end if;
	  else branch := branch_true; end if;
	  if hold_pc = '0' then
  	    if (branch = '1') then
              if (cond = BA) and (annul = '1') then annul_next := '1'; end if;
            else annul_next := annul; end if;
	    if r.d.inull = '1' then -- contention with JMPL
	      hold_pc := '1'; annul_current := '1'; annul_next := '0';
	    end if;
	  end if;
        end if;
      when FMT3 =>
        case op3 is
        when UMUL | SMUL | UMULCC | SMULCC =>
	  if true and (0 /= 0) then mulstart := '1'; end if;
	  if true and (0 = 0) then
            case r.d.cnt is
            when "00" =>
 	      cnt := "01"; hold_pc := '1'; pv := '0'; mulstart := '1';
            when "01" =>
 	      if mulo.nready = '1' then cnt := "00";
              else cnt := "01"; pv := '0'; hold_pc := '1'; end if;
            when others => null;
	    end case;
	  end if;
        when UDIV | SDIV | UDIVCC | SDIVCC =>
	  if true then
            case r.d.cnt is
            when "00" =>
 	      cnt := "01"; hold_pc := '1'; pv := '0';
	      divstart := '1';
            when "01" =>
 	      if divo.nready = '1' then cnt := "00"; 
              else cnt := "01"; pv := '0'; hold_pc := '1'; end if;
            when others => null;
	    end case;
	  end if;
        when TICC =>
	  if branch_true = '1' then ticc_exception := '1'; end if;
        when RETT =>
          rett_inst := '1'; --su := sregs.ps; 
        when JMPL =>
          de_jmpl := '1';
        when WRY =>
          if false then 
            if inst(29 downto 25) = "10011" then -- %ASR19
              case r.d.cnt is
              when "00" =>
                pv := '0'; cnt := "00"; hold_pc := '1';
                if r.x.ipend = '1' then cnt := "01"; end if;              
              when "01" =>
                cnt := "00";
              when others =>
              end case;
            end if;
          end if;
        when others => null;
        end case;
      when others =>  -- LDST 
        case r.d.cnt is
        when "00" =>
          if (op3(2) = '1') or (op3(1 downto 0) = "11") then -- ST/LDST/SWAP/LDD
 	    cnt := "01"; hold_pc := '1'; pv := '0';
          end if;
        when "01" =>
          if (op3(2 downto 0) = "111") or (op3(3 downto 0) = "1101") or
             ((false or FPEN) and ((op3(5) & op3(2 downto 0)) = "1110"))
	  then	-- LDD/STD/LDSTUB/SWAP
 	    cnt := "10"; pv := '0'; hold_pc := '1';
	  else
 	    cnt := "00";
          end if;
        when "10" =>
 	  cnt := "00";
        when others => null;
	end case;
      end case;
    end if;

    if ldlock = '1' then
      cnt := r.d.cnt; annul_next := '0'; pv := '1';
    end if;
    hold_pc := (hold_pc or ldlock) and not annul_all;

    if hold_pc = '1' then de_pc := r.d.pc; else de_pc := r.f.pc; end if;

    annul_current := (annul_current or ldlock or annul_all);
    ctrl_annul := r.d.annul or annul_all or annul_current;
    pv := pv and not ((r.d.inull and not hold_pc) or annul_all);
    jmpl_inst := de_jmpl and not annul_current;
    annul_next := (r.d.inull and not hold_pc) or annul_next or annul_all;
    if (annul_next = '1') or (rstn = '0') then
      cnt := (others => '0'); 
    end if;

    de_hold_pc := hold_pc; de_branch := branch; de_annul := annul_next;
    de_pv := pv; ctrl_pv := r.d.pv and 
	not ((r.d.annul and not r.d.pv) or annul_all or annul_current);
    inull := (not rstn) or r.d.inull or hold_pc or annul_all;

  end;

-- register write address generation

  procedure rd_gen(r : registers; inst : word; wreg, ld : out std_ulogic; 
	rdo : out std_logic_vector(4 downto 0)) is
  variable write_reg : std_ulogic;
  variable op : std_logic_vector(1 downto 0);
  variable op2 : std_logic_vector(2 downto 0);
  variable op3 : std_logic_vector(5 downto 0);
  variable rd  : std_logic_vector(4 downto 0);
  begin

    op    := inst(31 downto 30);
    op2   := inst(24 downto 22);
    op3   := inst(24 downto 19);

    write_reg := '0'; rd := inst(29 downto 25); ld := '0';

    case op is
    when CALL =>
        write_reg := '1'; rd := "01111";    -- CALL saves PC in r[15] (%o7)
    when FMT2 => 
        if (op2 = SETHI) then write_reg := '1'; end if;
    when FMT3 =>
        case op3 is
	when UMUL | SMUL | UMULCC | SMULCC => 
	  if true then
	    if (((mulo.nready = '1') and (r.d.cnt /= "00")) or (0 /= 0)) then
	      write_reg := '1'; 
	    end if;
	  else write_reg := '1'; end if;
	when UDIV | SDIV | UDIVCC | SDIVCC => 
	  if true then
	    if (divo.nready = '1') and (r.d.cnt /= "00") then
	      write_reg := '1'; 
	    end if;
	  else write_reg := '1'; end if;
        when RETT | WRPSR | WRY | WRWIM | WRTBR | TICC | FLUSH => null;
	when FPOP1 | FPOP2 => null;
	when CPOP1 | CPOP2 => null;
        when others => write_reg := '1';
        end case;
      when others =>   -- LDST
        ld := not op3(2);
        if (op3(2) = '0') and not ((false or FPEN) and (op3(5) = '1')) 
        then write_reg := '1'; end if;
        case op3 is
        when SWAP | SWAPA | LDSTUB | LDSTUBA =>
	  if r.d.cnt = "00" then write_reg := '1'; ld := '1'; end if;
        when others => null;
        end case;
        if r.d.cnt = "01" then
	  case op3 is
	  when LDD | LDDA | LDDC | LDDF => rd(0) := '1';
          when others =>
          end case;
      	end if;
    end case;

    if (rd = "00000") then write_reg := '0'; end if;
    wreg := write_reg; rdo := rd;
  end;

-- immediate data generation

  function imm_data (r : registers; insn : word) 
	return word is
  variable immediate_data, inst : word;
  begin
    immediate_data := (others => '0'); inst := insn;
    case inst(31 downto 30) is
    when FMT2 =>
      immediate_data := inst(21 downto 0) & "0000000000";
    when others =>	-- LDST
      immediate_data(31 downto 13) := (others => inst(12));
      immediate_data(12 downto 0) := inst(12 downto 0);
    end case;
    return(immediate_data);
  end;

-- read special registers
  function get_spr (r : registers) return word is
  variable spr : word;
  begin
    spr := (others => '0');
      case r.e.ctrl.inst(24 downto 19) is
      when RDPSR => spr(31 downto 5) := conv_std_logic_vector(15,4) &
        conv_std_logic_vector(3,4) & r.m.icc & "000000" & r.w.s.ec & r.w.s.ef & 
	r.w.s.pil & r.e.su & r.w.s.ps & r.e.et;
	spr(3-1 downto 0) := r.e.cwp;
      when RDTBR => spr(31 downto 4) := r.w.s.tba & r.w.s.tt;
      when RDWIM => spr(8-1 downto 0) := r.w.s.wim;
      when others =>
      end case;
    return(spr);
  end;

-- immediate data select

  function imm_select(inst : word) return boolean is
  variable imm : boolean;
  begin
    imm := false;
    case inst(31 downto 30) is
    when FMT2 =>
      case inst(24 downto 22) is
      when SETHI => imm := true;
      when others => 
      end case;
    when FMT3 =>
      case inst(24 downto 19) is
      when RDWIM | RDPSR | RDTBR => imm := true;
      when others => if (inst(13) = '1') then imm := true; end if;
      end case;
    when LDST => 
      if (inst(13) = '1') then imm := true; end if;
    when others => 
    end case;
    return(imm);
  end;

-- EXE operation

  procedure alu_op(r : in registers; iop1, iop2 : in word; me_icc : std_logic_vector(3 downto 0);
	my, ldbp : std_ulogic; aop1, aop2 : out word; aluop  : out std_logic_vector(2 downto 0);
	alusel : out std_logic_vector(1 downto 0); aluadd : out std_ulogic;
	shcnt : out std_logic_vector(4 downto 0); sari, shleft, ymsb, 
	mulins, divins, mulstep, macins, ldbp2, invop2 : out std_ulogic) is
  variable op : std_logic_vector(1 downto 0);
  variable op2 : std_logic_vector(2 downto 0);
  variable op3 : std_logic_vector(5 downto 0);
  variable rd  : std_logic_vector(4 downto 0);
  variable icc : std_logic_vector(3 downto 0);
  variable y0  : std_ulogic;
  begin

    op   := r.a.ctrl.inst(31 downto 30);
    op2  := r.a.ctrl.inst(24 downto 22);
    op3  := r.a.ctrl.inst(24 downto 19);
    aop1 := iop1; aop2 := iop2; ldbp2 := ldbp;
    aluop := EXE_NOP; alusel := EXE_RES_MISC; aluadd := '1'; 
    shcnt := iop2(4 downto 0); sari := '0'; shleft := '0'; invop2 := '0';
    ymsb := iop1(0); mulins := '0'; divins := '0'; mulstep := '0';
    macins := '0';

    if r.e.ctrl.wy = '1' then y0 := my;
    elsif r.m.ctrl.wy = '1' then y0 := r.m.y(0);
    elsif r.x.ctrl.wy = '1' then y0 := r.x.y(0);
    else y0 := r.w.s.y(0); end if;

    if r.e.ctrl.wicc = '1' then icc := me_icc;
    elsif r.m.ctrl.wicc = '1' then icc := r.m.icc;
    elsif r.x.ctrl.wicc = '1' then icc := r.x.icc;
    else icc := r.w.s.icc; end if;

    case op is
    when CALL =>
      aluop := EXE_LINK;
    when FMT2 =>
      case op2 is
      when SETHI => aluop := EXE_PASS2;
      when others =>
      end case;
    when FMT3 =>
      case op3 is
      when IADD | ADDX | ADDCC | ADDXCC | TADDCC | TADDCCTV | SAVE | RESTORE |
	   TICC | JMPL | RETT  => alusel := EXE_RES_ADD;
      when ISUB | SUBX | SUBCC | SUBXCC | TSUBCC | TSUBCCTV  => 
	alusel := EXE_RES_ADD; aluadd := '0'; aop2 := not iop2; invop2 := '1';
      when MULSCC => alusel := EXE_RES_ADD;
	aop1 := (icc(3) xor icc(1)) & iop1(31 downto 1);
	if y0 = '0' then aop2 := (others => '0'); ldbp2 := '0'; end if;
	mulstep := '1';
      when UMUL | UMULCC | SMUL | SMULCC => 
	if true then mulins := '1'; end if;
      when UMAC | SMAC => 
	if false then mulins := '1'; macins := '1'; end if;
      when UDIV | UDIVCC | SDIV | SDIVCC => 
	if true then 
	  aluop := EXE_DIV; alusel := EXE_RES_LOGIC; divins := '1';
        end if;
      when IAND | ANDCC => aluop := EXE_AND; alusel := EXE_RES_LOGIC;
      when ANDN | ANDNCC => aluop := EXE_ANDN; alusel := EXE_RES_LOGIC;
      when IOR | ORCC  => aluop := EXE_OR; alusel := EXE_RES_LOGIC;
      when ORN | ORNCC  => aluop := EXE_ORN; alusel := EXE_RES_LOGIC;
      when IXNOR | XNORCC  => aluop := EXE_XNOR; alusel := EXE_RES_LOGIC;
      when XORCC | IXOR | WRPSR | WRWIM | WRTBR | WRY  => 
	aluop := EXE_XOR; alusel := EXE_RES_LOGIC;
      when RDPSR | RDTBR | RDWIM => aluop := EXE_SPR;
      when RDY => aluop := EXE_RDY;
      when ISLL => aluop := EXE_SLL; alusel := EXE_RES_SHIFT; shleft := '1'; 
		   shcnt := not iop2(4 downto 0); invop2 := '1';
      when ISRL => aluop := EXE_SRL; alusel := EXE_RES_SHIFT; 
      when ISRA => aluop := EXE_SRA; alusel := EXE_RES_SHIFT; sari := iop1(31);
      when FPOP1 | FPOP2 =>
      when others =>
      end case;
    when others =>	-- LDST
      case r.a.ctrl.cnt is
      when "00" =>
        alusel := EXE_RES_ADD;
      when "01" =>
	case op3 is
	when LDD | LDDA | LDDC => alusel := EXE_RES_ADD;
	when LDDF => alusel := EXE_RES_ADD;
	when SWAP | SWAPA | LDSTUB | LDSTUBA => alusel := EXE_RES_ADD;
	when STF | STDF =>
	when others =>
          aluop := EXE_PASS1;
	  if op3(2) = '1' then 
	    if op3(1 downto 0) = "01" then aluop := EXE_STB;
	    elsif op3(1 downto 0) = "10" then aluop := EXE_STH; end if;
          end if;
        end case;
      when "10" =>
        aluop := EXE_PASS1;
        if op3(2) = '1' then  -- ST
          if (op3(3) and not op3(1))= '1' then aluop := EXE_ONES; end if; -- LDSTUB/A
        end if;
      when others =>
      end case;
    end case;
  end;

  function ra_inull_gen(r, v : registers) return std_ulogic is
  variable de_inull : std_ulogic;
  begin
    de_inull := '0';
    if ((v.e.jmpl or v.e.ctrl.rett) and not v.e.ctrl.annul and not (r.e.jmpl and not r.e.ctrl.annul)) = '1' then de_inull := '1'; end if;
    if ((v.a.jmpl or v.a.ctrl.rett) and not v.a.ctrl.annul and not (r.a.jmpl and not r.a.ctrl.annul)) = '1' then de_inull := '1'; end if;
    return(de_inull);
  end;

-- operand generation

  procedure op_mux(r : in registers; rfd, ed, md, xd, im : in word; 
	rsel : in std_logic_vector(2 downto 0); 
	ldbp : out std_ulogic; d : out word) is
  begin
    ldbp := '0';
    case rsel is
    when "000" => d := rfd;
    when "001" => d := ed;
    when "010" => d := md; if lddel = 1 then ldbp := r.m.ctrl.ld; end if;
    when "011" => d := xd;
    when "100" => d := im;
    when "101" => d := (others => '0');
    when "110" => d := r.w.result;
    when others => d := (others => '-');
    end case;
  end;

  procedure op_find(r : in registers; ldchkra : std_ulogic; ldchkex : std_ulogic;
	 rs1 : std_logic_vector(4 downto 0); ra : rfatype; im : boolean; rfe : out std_ulogic; 
	osel : out std_logic_vector(2 downto 0); ldcheck : std_ulogic) is
  begin
    rfe := '0';
    if im then osel := "100";
    elsif rs1 = "00000" then osel := "101";	-- %g0
    elsif ((r.a.ctrl.wreg and ldchkra) = '1') and (ra = r.a.ctrl.rd) then osel := "001";
    elsif ((r.e.ctrl.wreg and ldchkex) = '1') and (ra = r.e.ctrl.rd) then osel := "010";
    elsif r.m.ctrl.wreg = '1' and (ra = r.m.ctrl.rd) then osel := "011";
    elsif (irfwt = 0) and r.x.ctrl.wreg = '1' and (ra = r.x.ctrl.rd) then osel := "110";
    else  osel := "000"; rfe := ldcheck; end if;
  end;

-- generate carry-in for alu

  procedure cin_gen(r : registers; me_cin : in std_ulogic; cin : out std_ulogic) is
  variable op : std_logic_vector(1 downto 0);
  variable op3 : std_logic_vector(5 downto 0);
  variable ncin : std_ulogic;
  begin

    op := r.a.ctrl.inst(31 downto 30); op3 := r.a.ctrl.inst(24 downto 19);
    if r.e.ctrl.wicc = '1' then ncin := me_cin;
    else ncin := r.m.icc(0); end if;
    cin := '0';
    case op is
    when FMT3 =>
      case op3 is
      when ISUB | SUBCC | TSUBCC | TSUBCCTV => cin := '1';
      when ADDX | ADDXCC => cin := ncin; 
      when SUBX | SUBXCC => cin := not ncin; 
      when others => null;
      end case;
    when others => null;
    end case;
  end;

  procedure logic_op(r : registers; aluin1, aluin2, mey : word; 
	ymsb : std_ulogic; logicres, y : out word) is
  variable logicout : word;
  begin
    case r.e.aluop is
    when EXE_AND   => logicout := aluin1 and aluin2;
    when EXE_ANDN  => logicout := aluin1 and not aluin2;
    when EXE_OR    => logicout := aluin1 or aluin2;
    when EXE_ORN   => logicout := aluin1 or not aluin2;
    when EXE_XOR   => logicout := aluin1 xor aluin2;
    when EXE_XNOR  => logicout := aluin1 xor not aluin2;
    when EXE_DIV   => 
      if true then logicout := aluin2;
      else logicout := (others => '-'); end if;
    when others => logicout := (others => '-');
    end case;
    if (r.e.ctrl.wy and r.e.mulstep) = '1' then 
      y := ymsb & r.m.y(31 downto 1); 
    elsif r.e.ctrl.wy = '1' then y := logicout;
    elsif r.m.ctrl.wy = '1' then y := mey; 
    elsif false and (r.x.mac = '1') then y := mulo.result(63 downto 32);
    elsif r.x.ctrl.wy = '1' then y := r.x.y; 
    else y := r.w.s.y; end if;
    logicres := logicout;
  end;

  procedure misc_op(r : registers; wpr : watchpoint_registers; 
	aluin1, aluin2, ldata, mey : word; 
	mout, edata : out word) is
  variable miscout, bpdata, stdata : word;
  variable wpi : integer;
  begin
    wpi := 0; miscout := r.e.ctrl.pc(31 downto 2) & "00"; 
    edata := aluin1; bpdata := aluin1;
    if ((r.x.ctrl.wreg and r.x.ctrl.ld and not r.x.ctrl.annul) = '1') and
       (r.x.ctrl.rd = r.e.ctrl.rd) and (r.e.ctrl.inst(31 downto 30) = LDST) and
	(r.e.ctrl.cnt /= "10")
    then bpdata := ldata; end if;

    case r.e.aluop is
    when EXE_STB   => miscout := bpdata(7 downto 0) & bpdata(7 downto 0) &
			     bpdata(7 downto 0) & bpdata(7 downto 0);
		      edata := miscout;
    when EXE_STH   => miscout := bpdata(15 downto 0) & bpdata(15 downto 0);
		      edata := miscout;
    when EXE_PASS1 => miscout := bpdata; edata := miscout;
    when EXE_PASS2 => miscout := aluin2;
    when EXE_ONES  => miscout := (others => '1');
		      edata := miscout;
    when EXE_RDY  => 
      if true and (r.m.ctrl.wy = '1') then miscout := mey;
      else miscout := r.m.y; end if;
      if (NWP > 0) and (r.e.ctrl.inst(18 downto 17) = "11") then
 	wpi := conv_integer(r.e.ctrl.inst(16 downto 15));
 	if r.e.ctrl.inst(14) = '0' then miscout := wpr(wpi).addr & '0' & wpr(wpi).exec;
 	else miscout := wpr(wpi).mask & wpr(wpi).load & wpr(wpi).store; end if;
      end if;
      if (r.e.ctrl.inst(18 downto 17) = "10") and (r.e.ctrl.inst(14) = '1') then --%ASR17
        miscout := asr17_gen(r);
      end if;
      if false then
        if (r.e.ctrl.inst(18 downto 14) = "10010") then --%ASR18
          if ((r.m.mac = '1') and not false) or ((r.x.mac = '1') and false) then
            miscout := mulo.result(31 downto 0);	-- data forward of asr18
	  else miscout := r.w.s.asr18; end if;
        else
          if ((r.m.mac = '1') and not false) or ((r.x.mac = '1') and false) then
            miscout := mulo.result(63 downto 32);   -- data forward Y
	  end if;
        end if;
      end if;
    when EXE_SPR  => 
      miscout := get_spr(r);
    when others => null;
    end case;
    mout := miscout;
  end;

  procedure alu_select(r : registers; addout : std_logic_vector(32 downto 0);
	op1, op2 : word; shiftout, logicout, miscout : word; res : out word; 
	me_icc : std_logic_vector(3 downto 0);
	icco : out std_logic_vector(3 downto 0); divz : out std_ulogic) is
  variable op : std_logic_vector(1 downto 0);
  variable op3 : std_logic_vector(5 downto 0);
  variable icc : std_logic_vector(3 downto 0);
  variable aluresult : word;
  begin
    op   := r.e.ctrl.inst(31 downto 30); op3  := r.e.ctrl.inst(24 downto 19);
    icc := (others => '0');
    case r.e.alusel is
    when EXE_RES_ADD => 
      aluresult := addout(32 downto 1);
      if r.e.aluadd = '0' then
        icc(0) := ((not op1(31)) and not op2(31)) or 	-- Carry
		 (addout(32) and ((not op1(31)) or not op2(31)));
        icc(1) := (op1(31) and (op2(31)) and not addout(32)) or 	-- Overflow
                 (addout(32) and (not op1(31)) and not op2(31));
      else
        icc(0) := (op1(31) and op2(31)) or 	-- Carry
		 ((not addout(32)) and (op1(31) or op2(31)));
        icc(1) := (op1(31) and op2(31) and not addout(32)) or 	-- Overflow
		 (addout(32) and (not op1(31)) and (not op2(31)));
      end if;
      if notag = 0 then
        case op is 
        when FMT3 =>
          case op3 is
          when TADDCC | TADDCCTV =>
            icc(1) := op1(0) or op1(1) or op2(0) or op2(1) or icc(1);
          when TSUBCC | TSUBCCTV =>
            icc(1) := op1(0) or op1(1) or (not op2(0)) or (not op2(1)) or icc(1);
          when others => null;
          end case;
        when others => null;
        end case;
      end if;

      if aluresult = "00000000000000000000000000000000" then icc(2) := '1'; end if;
    when EXE_RES_SHIFT => aluresult := shiftout;
    when EXE_RES_LOGIC => aluresult := logicout;
      if aluresult = "00000000000000000000000000000000" then icc(2) := '1'; end if;
    when others => aluresult := miscout;
    end case;
    if r.e.jmpl = '1' then aluresult := r.e.ctrl.pc(31 downto 2) & "00"; end if;
    icc(3) := aluresult(31); divz := icc(2);
    if r.e.ctrl.wicc = '1' then
      if (op = FMT3) and (op3 = WRPSR) then icco := logicout(23 downto 20);
      else icco := icc; end if;
    elsif r.m.ctrl.wicc = '1' then icco := me_icc;
    elsif r.x.ctrl.wicc = '1' then icco := r.x.icc;
    else icco := r.w.s.icc; end if;
    res := aluresult;
  end;

  procedure dcache_gen(r, v : registers; dci : out dc_in_type; 
	link_pc, jump, force_a2, load : out std_ulogic) is
  variable op : std_logic_vector(1 downto 0);
  variable op3 : std_logic_vector(5 downto 0);
  variable su : std_ulogic;
  begin
    op := r.e.ctrl.inst(31 downto 30); op3 := r.e.ctrl.inst(24 downto 19);
    dci.signed := '0'; dci.lock := '0'; dci.dsuen := '0'; dci.size := SZWORD;
    if op = LDST then
    case op3 is
      when LDUB | LDUBA => dci.size := SZBYTE;
      when LDSTUB | LDSTUBA => dci.size := SZBYTE; dci.lock := '1'; 
      when LDUH | LDUHA => dci.size := SZHALF;
      when LDSB | LDSBA => dci.size := SZBYTE; dci.signed := '1';
      when LDSH | LDSHA => dci.size := SZHALF; dci.signed := '1';
      when LD | LDA | LDF | LDC => dci.size := SZWORD;
      when SWAP | SWAPA => dci.size := SZWORD; dci.lock := '1'; 
      when LDD | LDDA | LDDF | LDDC => dci.size := SZDBL;
      when STB | STBA => dci.size := SZBYTE;
      when STH | STHA => dci.size := SZHALF;
      when ST | STA | STF => dci.size := SZWORD;
      when ISTD | STDA => dci.size := SZDBL;
      when STDF | STDFQ => if FPEN then dci.size := SZDBL; end if;
      when STDC | STDCQ => if false then dci.size := SZDBL; end if;
      when others => dci.size := SZWORD; dci.lock := '0'; dci.signed := '0';
    end case;
    end if;
    
    link_pc := '0'; jump:= '0'; force_a2 := '0'; load := '0';
    dci.write := '0'; dci.enaddr := '0'; dci.read := not op3(2);

-- load/store control decoding

    if (r.e.ctrl.annul = '0') then
      case op is
      when CALL => link_pc := '1';
      when FMT3 =>
        case op3 is
        when JMPL => jump := '1'; link_pc := '1'; 
        when RETT => jump := '1';
        when others => null;
        end case;
      when LDST =>
          case r.e.ctrl.cnt is
	  when "00" =>
            dci.read := op3(3) or not op3(2);	-- LD/LDST/SWAP
            load := op3(3) or not op3(2);
	    dci.enaddr := '1';
          when "01" =>
            force_a2 := not op3(2);	-- LDD
            load := not op3(2); dci.enaddr := not op3(2);
            if op3(3 downto 2) = "01" then		-- ST/STD
	      dci.write := '1';
            end if;
            if op3(3 downto 2) = "11" then		-- LDST/SWAP
	      dci.enaddr := '1';
            end if;
          when "10" => 					-- STD/LDST/SWAP
            dci.write := '1';
          when others => null;
	  end case;
	if (r.e.ctrl.trap or (v.x.ctrl.trap and not v.x.ctrl.annul)) = '1' then
	  dci.enaddr := '0';
	end if;
      when others => null;
      end case;
    end if;

    if ((r.x.ctrl.rett and not r.x.ctrl.annul) = '1') then su := r.w.s.ps;
    else su := r.w.s.s; end if;
    if su = '1' then dci.asi := "00001011"; else dci.asi := "00001010"; end if;
    if (op3(4) = '1') and ((op3(5) = '0') or not false) then
      dci.asi := r.e.ctrl.inst(12 downto 5);
    end if;

  end;

  procedure fpstdata(r : in registers; edata, eres : in word; fpstdata : in std_logic_vector(31 downto 0);
                       edata2, eres2 : out word) is
    variable op : std_logic_vector(1 downto 0);
    variable op3 : std_logic_vector(5 downto 0);
  begin
    edata2 := edata; eres2 := eres;
    op := r.e.ctrl.inst(31 downto 30); op3 := r.e.ctrl.inst(24 downto 19);
    if FPEN then
      if FPEN and (op = LDST) and  ((op3(5 downto 4) & op3(2)) = "101") and (r.e.ctrl.cnt /= "00") then
        edata2 := fpstdata; eres2 := fpstdata;
      end if;
    end if;
  end;
  
  function ld_align(data : dcdtype; set : std_logic_vector(0 downto 0);
	size, laddr : std_logic_vector(1 downto 0); signed : std_ulogic) return word is
  variable align_data, rdata : word;
  begin
    align_data := data(conv_integer(set)); rdata := (others => '0');
    case size is
    when "00" => 			-- byte read
      case laddr is
      when "00" => 
	rdata(7 downto 0) := align_data(31 downto 24);
	if signed = '1' then rdata(31 downto 8) := (others => align_data(31)); end if;
      when "01" => 
	rdata(7 downto 0) := align_data(23 downto 16);
	if signed = '1' then rdata(31 downto 8) := (others => align_data(23)); end if;
      when "10" => 
	rdata(7 downto 0) := align_data(15 downto 8);
	if signed = '1' then rdata(31 downto 8) := (others => align_data(15)); end if;
      when others => 
	rdata(7 downto 0) := align_data(7 downto 0);
	if signed = '1' then rdata(31 downto 8) := (others => align_data(7)); end if;
      end case;
    when "01" => 			-- half-word read
      if  laddr(1) = '1' then 
	rdata(15 downto 0) := align_data(15 downto 0);
	if signed = '1' then rdata(31 downto 15) := (others => align_data(15)); end if;
      else
	rdata(15 downto 0) := align_data(31 downto 16);
	if signed = '1' then rdata(31 downto 15) := (others => align_data(31)); end if;
      end if;
    when others => 			-- single and double word read
      rdata := align_data;
    end case;
    return(rdata);
  end;

  procedure mem_trap(r : registers; wpr : watchpoint_registers;
                     annul, holdn : in std_ulogic;
                     trapout, iflush, nullify, werrout : out std_ulogic;
                     tt : out std_logic_vector(5 downto 0)) is
  variable cwp   : std_logic_vector(3-1 downto 0);
  variable cwpx  : std_logic_vector(5 downto 3);
  variable op : std_logic_vector(1 downto 0);
  variable op2 : std_logic_vector(2 downto 0);
  variable op3 : std_logic_vector(5 downto 0);
  variable nalign_d : std_ulogic;
  variable trap, werr : std_ulogic;
  begin
    op := r.m.ctrl.inst(31 downto 30); op2  := r.m.ctrl.inst(24 downto 22);
    op3 := r.m.ctrl.inst(24 downto 19);
    cwpx := r.m.result(5 downto 3); cwpx(5) := '0';
    iflush := '0'; trap := r.m.ctrl.trap; nullify := annul;
    tt := r.m.ctrl.tt; werr := (dco.werr or r.m.werr) and not r.w.s.dwt;
    nalign_d := r.m.nalign or r.m.result(2); 
    if ((annul or trap) /= '1') and (r.m.ctrl.pv = '1') then
      if (werr and holdn) = '1' then
	trap := '1'; tt := TT_DSEX; werr := '0';
        if op = LDST then nullify := '1'; end if;
      end if;
    end if;
    if ((annul or trap) /= '1') then      
      case op is
      when FMT2 =>
        case op2 is
        when FBFCC => 
          if FPEN and (fpo.exc = '1') then trap := '1'; tt := TT_FPEXC; end if;
        when CBCCC =>
    	  if false and (cpo.exc = '1') then trap := '1'; tt := TT_CPEXC; end if;
        when others => null;
        end case;
      when FMT3 =>
        case op3 is
	when WRPSR =>
	  if (orv(cwpx) = '1') then trap := '1'; tt := TT_IINST; end if;
	when UDIV | SDIV | UDIVCC | SDIVCC =>
    	  if true then 
	    if r.m.divz = '1' then trap := '1'; tt := TT_DIV; end if;
          end if;
	when JMPL | RETT =>
	  if r.m.nalign = '1' then trap := '1'; tt := TT_UNALA; end if;
        when TADDCCTV | TSUBCCTV =>
	  if (notag = 0) and (r.m.icc(1) = '1') then
	    trap := '1'; tt := TT_TAG;
	  end if;
	when FLUSH => iflush := '1';
	when FPOP1 | FPOP2 =>
          if FPEN and (fpo.exc = '1') then trap := '1'; tt := TT_FPEXC; end if;
	when CPOP1 | CPOP2 =>
    	  if false and (cpo.exc = '1') then trap := '1'; tt := TT_CPEXC; end if;
        when others => null;
        end case;
      when LDST =>
        if r.m.ctrl.cnt = "00" then
          case op3 is
            when LDDF | STDF | STDFQ =>
	    if FPEN then
	      if nalign_d = '1' then
	        trap := '1'; tt := TT_UNALA; nullify := '1';
              elsif (fpo.exc and r.m.ctrl.pv) = '1' 
              then trap := '1'; tt := TT_FPEXC; nullify := '1'; end if;
	    end if;
	  when LDDC | STDC | STDCQ =>
	    if false then
	      if nalign_d = '1' then
	        trap := '1'; tt := TT_UNALA; nullify := '1';
    	      elsif ((cpo.exc and r.m.ctrl.pv) = '1') 
    	      then trap := '1'; tt := TT_CPEXC; nullify := '1'; end if;
	    end if;
	  when LDD | ISTD | LDDA | STDA =>
	    if r.m.result(2 downto 0) /= "000" then
	      trap := '1'; tt := TT_UNALA; nullify := '1';
	    end if;
 	  when LDF | LDFSR | STFSR | STF =>
	    if FPEN and (r.m.nalign = '1') then
	      trap := '1'; tt := TT_UNALA; nullify := '1';
            elsif FPEN and ((fpo.exc and r.m.ctrl.pv) = '1')
            then trap := '1'; tt := TT_FPEXC; nullify := '1'; end if;
 	  when LDC | LDCSR | STCSR | STC =>
	    if false and (r.m.nalign = '1') then 
	      trap := '1'; tt := TT_UNALA; nullify := '1';
    	    elsif false and ((cpo.exc and r.m.ctrl.pv) = '1') 
    	    then trap := '1'; tt := TT_CPEXC; nullify := '1'; end if;
 	  when LD | LDA | ST | STA | SWAP | SWAPA =>
	    if r.m.result(1 downto 0) /= "00" then
	      trap := '1'; tt := TT_UNALA; nullify := '1';
	    end if;
          when LDUH | LDUHA | LDSH | LDSHA | STH | STHA =>
	    if r.m.result(0) /= '0' then
	      trap := '1'; tt := TT_UNALA; nullify := '1';
	    end if;
          when others => null;
          end case;
          for i in 1 to NWP loop
            if ((((wpr(i-1).load and not op3(2)) or (wpr(i-1).store and op3(2))) = '1') and
                (((wpr(i-1).addr xor r.m.result(31 downto 2)) and wpr(i-1).mask) = "000000000000000000000000000000"))
            then trap := '1'; tt := TT_WATCH; nullify := '1'; end if;
          end loop;
	end if;
      when others => null;
      end case;
    end if;
    if (rstn = '0') or (r.x.rstate = dsu2) then werr := '0'; end if;
    trapout := trap; werrout := werr;
  end;

  procedure irq_trap(r       : in registers;
                     ir      : in irestart_register;
                     irl     : in std_logic_vector(3 downto 0);
                     annul   : in std_ulogic;
                     pv      : in std_ulogic;
                     trap    : in std_ulogic;
                     tt      : in std_logic_vector(5 downto 0);
                     nullify : in std_ulogic;
                     irqen   : out std_ulogic;
                     irqen2  : out std_ulogic;
                     nullify2 : out std_ulogic;
                     trap2, ipend  : out std_ulogic;
                     tt2      : out std_logic_vector(5 downto 0)) is
    variable op : std_logic_vector(1 downto 0);
    variable op3 : std_logic_vector(5 downto 0);
    variable pend : std_ulogic;
  begin
    nullify2 := nullify; trap2 := trap; tt2 := tt; 
    op := r.m.ctrl.inst(31 downto 30); op3 := r.m.ctrl.inst(24 downto 19);
    irqen := '1'; irqen2 := r.m.irqen;

    if (annul or trap) = '0' then
      if ((op = FMT3) and (op3 = WRPSR)) then irqen := '0'; end if;    
    end if;

    if (irl = "1111") or (irl > r.w.s.pil) then
      pend := r.m.irqen and r.m.irqen2 and r.w.s.et and not ir.pwd;
    else pend := '0'; end if;
    ipend := pend;

    if ((not annul) and pv and (not trap) and pend) = '1' then
      trap2 := '1'; tt2 := "01" & irl;
      if op = LDST then nullify2 := '1'; end if;
    end if;
  end;

  procedure irq_intack(r : in registers; holdn : in std_ulogic; intack: out std_ulogic) is 
  begin
    intack := '0';
    if r.x.rstate = trap then 
      if r.w.s.tt(7 downto 4) = "0001" then intack := '1'; end if;
    end if;
  end;
  
-- write special registers

  procedure sp_write (r : registers; wpr : watchpoint_registers;
        s : out special_register_type; vwpr : out watchpoint_registers) is
  variable op : std_logic_vector(1 downto 0);
  variable op2 : std_logic_vector(2 downto 0);
  variable op3 : std_logic_vector(5 downto 0);
  variable rd  : std_logic_vector(4 downto 0);
  variable i   : integer range 0 to 3;
  begin

    op  := r.x.ctrl.inst(31 downto 30);
    op2 := r.x.ctrl.inst(24 downto 22);
    op3 := r.x.ctrl.inst(24 downto 19);
    s   := r.w.s;
    rd  := r.x.ctrl.inst(29 downto 25);
    vwpr := wpr;
    
      case op is
      when FMT3 =>
        case op3 is
        when WRY =>
          if rd = "00000" then
            s.y := r.x.result;
          elsif false and (rd = "10010") then
	    s.asr18 := r.x.result;
          elsif (rd = "10001") then
	    s.dwt := r.x.result(14);
            if (svt = 1) then s.svt := r.x.result(13); end if;
          elsif rd(4 downto 3) = "11" then -- %ASR24 - %ASR31
	    case rd(2 downto 0) is
	    when "000" => 
              vwpr(0).addr := r.x.result(31 downto 2);
              vwpr(0).exec := r.x.result(0); 
	    when "001" => 
              vwpr(0).mask := r.x.result(31 downto 2);
              vwpr(0).load := r.x.result(1);
              vwpr(0).store := r.x.result(0);              
	    when "010" => 
              vwpr(1).addr := r.x.result(31 downto 2);
              vwpr(1).exec := r.x.result(0); 
	    when "011" => 
              vwpr(1).mask := r.x.result(31 downto 2);
              vwpr(1).load := r.x.result(1);
              vwpr(1).store := r.x.result(0);              
	    when "100" => 
              vwpr(2).addr := r.x.result(31 downto 2);
              vwpr(2).exec := r.x.result(0); 
	    when "101" => 
              vwpr(2).mask := r.x.result(31 downto 2);
              vwpr(2).load := r.x.result(1);
              vwpr(2).store := r.x.result(0);              
	    when "110" => 
              vwpr(3).addr := r.x.result(31 downto 2);
              vwpr(3).exec := r.x.result(0); 
	    when others =>   -- "111"
              vwpr(3).mask := r.x.result(31 downto 2);
              vwpr(3).load := r.x.result(1);
              vwpr(3).store := r.x.result(0);              
            end case;
          end if;
        when WRPSR =>
          s.cwp := r.x.result(3-1 downto 0);
          s.icc := r.x.result(23 downto 20);
          s.ec  := r.x.result(13);
          if FPEN then s.ef  := r.x.result(12); end if;
          s.pil := r.x.result(11 downto 8);
          s.s   := r.x.result(7);
          s.ps  := r.x.result(6);
          s.et  := r.x.result(5);
        when WRWIM =>
          s.wim := r.x.result(8-1 downto 0);
        when WRTBR =>
          s.tba := r.x.result(31 downto 12);
        when SAVE =>
          if (not true) and (r.w.s.cwp = "000") then s.cwp := "111";
          else s.cwp := r.w.s.cwp - 1 ; end if;
        when RESTORE =>
          if (not true) and (r.w.s.cwp = "111") then s.cwp := "000";
          else s.cwp := r.w.s.cwp + 1; end if;
        when RETT =>
          if (not true) and (r.w.s.cwp = "111") then s.cwp := "000";
          else s.cwp := r.w.s.cwp + 1; end if;
          s.s := r.w.s.ps;
          s.et := '1';
        when others => null;
        end case;
      when others => null;
      end case;
      if r.x.ctrl.wicc = '1' then s.icc := r.x.icc; end if;
      if r.x.ctrl.wy = '1' then s.y := r.x.y; end if;
      if false and (r.x.mac = '1') then 
        s.asr18 := mulo.result(31 downto 0);
	s.y := mulo.result(63 downto 32);
      end if;
  end;

  function npc_find (r : registers) return std_logic_vector is
  variable npc : std_logic_vector(2 downto 0);
  begin
    npc := "011";
    if r.m.ctrl.pv = '1' then npc := "000";
    elsif r.e.ctrl.pv = '1' then npc := "001";
    elsif r.a.ctrl.pv = '1' then npc := "010";
    elsif r.d.pv = '1' then npc := "011";
    elsif 2 /= 0 then npc := "100"; end if;
    return(npc);
  end;

  function npc_gen (r : registers) return word is
  variable npc : std_logic_vector(31 downto 0);
  begin
    npc :=  r.a.ctrl.pc(31 downto 2) & "00";
    case r.x.npc is
    when "000" => npc(31 downto 2) := r.x.ctrl.pc(31 downto 2);
    when "001" => npc(31 downto 2) := r.m.ctrl.pc(31 downto 2);
    when "010" => npc(31 downto 2) := r.e.ctrl.pc(31 downto 2);
    when "011" => npc(31 downto 2) := r.a.ctrl.pc(31 downto 2);
    when others => 
	if 2 /= 0 then npc(31 downto 2) := r.d.pc(31 downto 2); end if;
    end case;
    return(npc);
  end;

  procedure mul_res(r : registers; asr18in : word; result, y, asr18 : out word; 
	  icc : out std_logic_vector(3 downto 0)) is
  variable op  : std_logic_vector(1 downto 0);
  variable op3 : std_logic_vector(5 downto 0);
  begin
    op    := r.m.ctrl.inst(31 downto 30); op3   := r.m.ctrl.inst(24 downto 19);
    result := r.m.result; y := r.m.y; icc := r.m.icc; asr18 := asr18in;
    case op is
    when FMT3 =>
      case op3 is
      when UMUL | SMUL =>
    	if true then 
	  result := mulo.result(31 downto 0);
          y := mulo.result(63 downto 32);
        end if;
      when UMULCC | SMULCC =>
    	if true then 
          result := mulo.result(31 downto 0); icc := mulo.icc;
          y := mulo.result(63 downto 32);
        end if;
      when UMAC | SMAC =>
	if false and not false then
	  result := mulo.result(31 downto 0);
	  asr18  := mulo.result(31 downto 0);
          y := mulo.result(63 downto 32);
	end if;
      when UDIV | SDIV =>
    	if true then 
          result := divo.result(31 downto 0);
        end if;
      when UDIVCC | SDIVCC =>
    	if true then 
          result := divo.result(31 downto 0); icc := divo.icc;
        end if;
      when others => null;
      end case;
    when others => null;
    end case;
  end;

  function powerdwn(r : registers; trap : std_ulogic; rp : pwd_register_type) return std_ulogic is
    variable op : std_logic_vector(1 downto 0);
    variable op3 : std_logic_vector(5 downto 0);
    variable rd  : std_logic_vector(4 downto 0);
    variable pd  : std_ulogic;
  begin
    op := r.x.ctrl.inst(31 downto 30);
    op3 := r.x.ctrl.inst(24 downto 19);
    rd  := r.x.ctrl.inst(29 downto 25);    
    pd := '0';
    if (not (r.x.ctrl.annul or trap) and r.x.ctrl.pv) = '1' then
      if ((op = FMT3) and (op3 = WRY) and (rd = "10011")) then pd := '1'; end if;
      pd := pd or rp.pwd;
    end if;
    return(pd);
  end;
  
  signal dummy : std_ulogic;
  signal cpu_index : std_logic_vector(3 downto 0);
  signal disasen : std_ulogic;

-- Signals used for tracking if a handler fired and which one
signal dfp_trap_vector : std_logic_vector(3129 downto 0);
signal or_reduce_1 : std_logic;
signal dfp_delay_start : integer range 0 to 15;
signal dfp_trap_mem : std_logic_vector(dfp_trap_vector'left downto dfp_trap_vector'right);
signal handlerTrap : std_ulogic;

-- Signals that serve as shadow signals for variables used in the pairs
signal V_A_ET_shadow : STD_ULOGIC;
signal EX_ADD_RES32DOWNTO34DOWNTO3_shadow : STD_LOGIC_VECTOR(4 downto 3);
signal ICNT_shadow : STD_ULOGIC;
signal EX_OP1_shadow : WORD;
signal V_M_CTRL_PC_shadow : PCTYPE;
signal V_E_CTRL_PC3DOWNTO2_shadow : std_logic_vector(3 downto 2);
signal DE_REN1_shadow : STD_ULOGIC;
signal DE_INST_shadow : WORD;
signal V_A_CTRL_CNT_shadow : OP_TYPE;
signal V_F_PC3DOWNTO2_shadow : std_logic_vector(3 downto 2);
signal V_W_S_TT_shadow : STD_LOGIC_VECTOR(7 downto 0);
signal V_X_RESULT6DOWNTO0_shadow : std_logic_vector(6 downto 0);
signal EX_JUMP_ADDRESS3DOWNTO2_shadow : std_logic_vector(3 downto 2);
signal V_E_ALUCIN_shadow : STD_ULOGIC;
signal V_D_PC3DOWNTO2_shadow : std_logic_vector(3 downto 2);
signal V_A_CTRL_PV_shadow : STD_ULOGIC;
signal V_E_CTRL_shadow : PIPELINE_CTRL_TYPE;
signal V_M_CTRL_shadow : PIPELINE_CTRL_TYPE;
signal V_M_RESULT1DOWNTO0_shadow : std_logic_vector(1 downto 0);
signal EX_SHCNT_shadow : ASI_TYPE;
signal V_M_DCI_SIZE_shadow : OP_TYPE;
signal V_X_CTRL_ANNUL_shadow : STD_ULOGIC;
signal V_X_MEXC_shadow : STD_ULOGIC;
signal TBUFCNTX_shadow : STD_LOGIC_VECTOR(6 downto 0);
signal V_A_CTRL_WY_shadow : STD_ULOGIC;
signal NPC_shadow : PCTYPE;
signal V_M_CTRL_TT3DOWNTO0_shadow : std_logic_vector(3 downto 0);
signal V_A_MULSTART_shadow : STD_ULOGIC;
signal XC_VECTT3DOWNTO0_shadow : STD_LOGIC_VECTOR(3 downto 0);
signal V_E_CTRL_TT_shadow : OP3_TYPE;
signal DSIGN_shadow : STD_ULOGIC;
signal V_E_CTRL_ANNUL_shadow : STD_ULOGIC;
signal EX_JUMP_ADDRESS_shadow : PCTYPE;
signal V_A_CTRL_PC31DOWNTO12_shadow : std_logic_vector(31 downto 12);
signal V_A_RFE1_shadow : STD_ULOGIC;
signal V_W_WA_shadow : RFATYPE;
signal V_X_ANNUL_ALL_shadow : STD_ULOGIC;
signal EX_YMSB_shadow : STD_ULOGIC;
signal EX_ADD_RES_shadow : STD_LOGIC_VECTOR(32 downto 0);
signal VIR_ADDR_shadow : PCTYPE;
signal EX_JUMP_ADDRESS31DOWNTO12_shadow : std_logic_vector(31 downto 12);
signal V_W_S_CWP_shadow : CWPTYPE;
signal V_D_INST0_shadow : std_logic_vector(31 downto 0);
signal V_A_CTRL_ANNUL_shadow : STD_ULOGIC;
signal V_X_DATA1_shadow : std_logic_vector(31 downto 0);
signal VP_PWD_shadow : STD_ULOGIC;
signal V_M_CTRL_RD6DOWNTO0_shadow : std_logic_vector(6 downto 0);
signal V_X_DATA00_shadow : STD_LOGIC;
signal V_M_CTRL_RETT_shadow : STD_ULOGIC;
signal V_X_CTRL_RETT_shadow : STD_ULOGIC;
signal V_X_CTRL_PC31DOWNTO12_shadow : std_logic_vector(31 downto 12);
signal V_W_S_PS_shadow : STD_ULOGIC;
signal V_X_CTRL_TT_shadow : OP3_TYPE;
signal V_D_STEP_shadow : STD_ULOGIC;
signal V_X_CTRL_WICC_shadow : STD_ULOGIC;
signal VIR_ADDR31DOWNTO2_shadow : std_logic_vector(31 downto 2);
signal V_M_CTRL_RD7DOWNTO0_shadow : std_logic_vector(7 downto 0);
signal V_X_RESULT_shadow : WORD;
signal V_D_CNT_shadow : OP_TYPE;
signal XC_VECTT_shadow : STD_LOGIC_VECTOR(7 downto 0);
signal EX_ADD_RES32DOWNTO3_shadow : STD_LOGIC_VECTOR(32 downto 3);
signal V_W_S_EF_shadow : STD_ULOGIC;
signal V_A_CTRL_PC31DOWNTO2_shadow : std_logic_vector(31 downto 2);
signal V_X_DATA04DOWNTO0_shadow : std_logic_vector(4 downto 0);
signal V_X_DCI_SIGNED_shadow : STD_ULOGIC;
signal V_M_NALIGN_shadow : STD_ULOGIC;
signal XC_WREG_shadow : STD_ULOGIC;
signal V_A_RFA2_shadow : RFATYPE;
signal V_E_CTRL_PC31DOWNTO12_shadow : std_logic_vector(31 downto 12);
signal EX_ADD_RES32DOWNTO332DOWNTO13_shadow : STD_LOGIC_VECTOR(32 downto 13);
signal EX_OP231_shadow : STD_LOGIC;
signal XC_TRAP_ADDRESS31DOWNTO4_shadow : std_logic_vector(31 downto 4);
signal V_X_ICC_shadow : STD_LOGIC_VECTOR(3 downto 0);
signal V_A_SU_shadow : STD_ULOGIC;
signal V_E_OP2_shadow : WORD;
signal EX_FORCE_A2_shadow : STD_ULOGIC;
signal V_E_CTRL_PC31DOWNTO2_shadow : std_logic_vector(31 downto 2);
signal V_E_CTRL_PC31DOWNTO4_shadow : std_logic_vector(31 downto 4);
signal V_E_OP131_shadow : STD_LOGIC;
signal V_X_DCI_shadow : DC_IN_TYPE;
signal V_E_CTRL_WICC_shadow : STD_ULOGIC;
signal EX_OP13_shadow : STD_LOGIC;
signal V_F_PC31DOWNTO12_shadow : std_logic_vector(31 downto 12);
signal V_E_CTRL_INST_shadow : WORD;
signal V_E_CTRL_LD_shadow : STD_ULOGIC;
signal V_M_SU_shadow : STD_ULOGIC;
signal V_E_SARI_shadow : STD_ULOGIC;
signal V_E_ET_shadow : STD_ULOGIC;
signal V_M_CTRL_PV_shadow : STD_ULOGIC;
signal VDSU_CRDY2_shadow : STD_LOGIC;
signal MUL_OP2_shadow : WORD;
signal XC_EXCEPTION_shadow : STD_ULOGIC;
signal V_E_OP1_shadow : WORD;
signal VP_ERROR_shadow : STD_ULOGIC;
signal V_M_DCI_SIGNED_shadow : STD_ULOGIC;
signal V_D_PC31DOWNTO12_shadow : std_logic_vector(31 downto 12);
signal MUL_OP231_shadow : STD_LOGIC;
signal XC_TRAP_ADDRESS31DOWNTO2_shadow : std_logic_vector(31 downto 2);
signal V_M_CTRL_PC3DOWNTO2_shadow : std_logic_vector(3 downto 2);
signal V_M_DCI_shadow : DC_IN_TYPE;
signal EX_OP23_shadow : STD_LOGIC;
signal V_X_CTRL_RD6DOWNTO0_shadow : std_logic_vector(6 downto 0);
signal V_X_CTRL_TRAP_shadow : STD_ULOGIC;
signal V_A_DIVSTART_shadow : STD_ULOGIC;
signal V_X_RESULT6DOWNTO03DOWNTO0_shadow : std_logic_vector(3 downto 0);
signal VDSU_TT_shadow : STD_LOGIC_VECTOR(7 downto 0);
signal EX_ADD_RES32DOWNTO332DOWNTO5_shadow : STD_LOGIC_VECTOR(32 downto 5);
signal V_X_CTRL_CNT_shadow : OP_TYPE;
signal V_E_YMSB_shadow : STD_ULOGIC;
signal EX_ADD_RES32DOWNTO330DOWNTO11_shadow : STD_LOGIC_VECTOR(30 downto 11);
signal V_A_RFE2_shadow : STD_ULOGIC;
signal V_E_OP13_shadow : STD_LOGIC;
signal V_A_CWP_shadow : CWPTYPE;
signal ME_SIZE_shadow : OP_TYPE;
signal V_X_MAC_shadow : STD_ULOGIC;
signal V_M_CTRL_INST_shadow : WORD;
signal VIR_ADDR31DOWNTO4_shadow : std_logic_vector(31 downto 4);
signal V_A_CTRL_INST20_shadow : STD_LOGIC;
signal DE_REN2_shadow : STD_ULOGIC;
signal V_E_CTRL_PV_shadow : STD_ULOGIC;
signal V_E_MAC_shadow : STD_ULOGIC;
signal V_X_CTRL_TT3DOWNTO0_shadow : std_logic_vector(3 downto 0);
signal EX_ADD_RES3_shadow : STD_LOGIC;
signal V_X_CTRL_INST_shadow : WORD;
signal V_M_CTRL_PC31DOWNTO2_shadow : std_logic_vector(31 downto 2);
signal V_W_S_ET_shadow : STD_ULOGIC;
signal V_M_CTRL_CNT_shadow : OP_TYPE;
signal V_M_CTRL_ANNUL_shadow : STD_ULOGIC;
signal DE_INST19_shadow : STD_LOGIC;
signal XC_HALT_shadow : STD_ULOGIC;
signal V_E_OP231_shadow : STD_LOGIC;
signal V_A_CTRL_PC3DOWNTO2_shadow : std_logic_vector(3 downto 2);
signal VIR_ADDR31DOWNTO12_shadow : std_logic_vector(31 downto 12);
signal V_M_CTRL_WICC_shadow : STD_ULOGIC;
signal V_M_CTRL_WREG_shadow : STD_ULOGIC;
signal V_W_S_S_shadow : STD_ULOGIC;
signal V_F_PC31DOWNTO2_shadow : std_logic_vector(31 downto 2);
signal V_E_CWP_shadow : CWPTYPE;
signal V_A_STEP_shadow : STD_ULOGIC;
signal V_A_CTRL_TT3DOWNTO0_shadow : std_logic_vector(3 downto 0);
signal V_A_CTRL_TRAP_shadow : STD_ULOGIC;
signal NPC31DOWNTO2_shadow : std_logic_vector(31 downto 2);
signal V_M_CTRL_TRAP_shadow : STD_ULOGIC;
signal V_D_PC31DOWNTO4_shadow : std_logic_vector(31 downto 4);
signal V_X_INTACK_shadow : STD_ULOGIC;
signal SIDLE_shadow : STD_ULOGIC;
signal V_A_CTRL_RETT_shadow : STD_ULOGIC;
signal V_X_DATA03_shadow : STD_LOGIC;
signal V_A_CTRL_INST19_shadow : STD_LOGIC;
signal V_W_S_SVT_shadow : STD_ULOGIC;
signal V_A_CTRL_PC31DOWNTO4_shadow : std_logic_vector(31 downto 4);
signal V_X_LADDR_shadow : OP_TYPE;
signal V_W_S_DWT_shadow : STD_ULOGIC;
signal EX_JUMP_ADDRESS31DOWNTO2_shadow : std_logic_vector(31 downto 2);
signal V_W_S_TBA_shadow : STD_LOGIC_VECTOR(19 downto 0);
signal XC_WADDR6DOWNTO0_shadow : STD_LOGIC_VECTOR(6 downto 0);
signal V_M_MUL_shadow : STD_ULOGIC;
signal V_E_SU_shadow : STD_ULOGIC;
signal V_M_Y31_shadow : STD_LOGIC;
signal V_E_OP23_shadow : STD_LOGIC;
signal V_M_CTRL_PC31DOWNTO4_shadow : std_logic_vector(31 downto 4);
signal DE_RADDR17DOWNTO0_shadow : STD_LOGIC_VECTOR(7 downto 0);
signal V_X_CTRL_PC31DOWNTO2_shadow : std_logic_vector(31 downto 2);
signal V_E_CTRL_TRAP_shadow : STD_ULOGIC;
signal V_X_DEBUG_shadow : STD_ULOGIC;
signal V_M_DCI_LOCK_shadow : STD_ULOGIC;
signal V_X_CTRL_PC3DOWNTO2_shadow : std_logic_vector(3 downto 2);
signal V_X_CTRL_WREG_shadow : STD_ULOGIC;
signal V_E_CTRL_INST24_shadow : STD_LOGIC;
signal V_D_MEXC_shadow : STD_ULOGIC;
signal V_W_RESULT_shadow : WORD;
signal VFPI_DBG_ENABLE_shadow : STD_ULOGIC;
signal EX_OP131_shadow : STD_LOGIC;
signal V_D_INST1_shadow : std_logic_vector(31 downto 0);
signal V_W_EXCEPT_shadow : STD_ULOGIC;
signal V_E_CTRL_TT3DOWNTO0_shadow : std_logic_vector(3 downto 0);
signal ME_LADDR_shadow : OP_TYPE;
signal V_X_CTRL_PC31DOWNTO4_shadow : std_logic_vector(31 downto 4);
signal V_E_CTRL_RETT_shadow : STD_ULOGIC;
signal XC_WADDR7DOWNTO0_shadow : STD_LOGIC_VECTOR(7 downto 0);
signal V_X_CTRL_PV_shadow : STD_ULOGIC;
signal V_E_CTRL_RD6DOWNTO0_shadow : std_logic_vector(6 downto 0);
signal V_M_MAC_shadow : STD_ULOGIC;
signal V_D_SET_shadow : STD_LOGIC_VECTOR(0 downto 0);
signal VIR_ADDR3DOWNTO2_shadow : std_logic_vector(3 downto 2);
signal V_D_CWP_shadow : CWPTYPE;
signal DE_INST20_shadow : STD_LOGIC;
signal V_D_ANNUL_shadow : STD_ULOGIC;
signal EX_OP2_shadow : WORD;
signal EX_SARI_shadow : STD_ULOGIC;
signal V_D_PC31DOWNTO2_shadow : std_logic_vector(31 downto 2);
signal V_X_DCI_SIZE_shadow : OP_TYPE;
signal V_M_Y_shadow : WORD;
signal V_X_CTRL_PC_shadow : PCTYPE;
signal V_X_SET_shadow : STD_LOGIC_VECTOR(0 downto 0);
signal V_A_CTRL_PC_shadow : PCTYPE;
signal V_A_JMPL_shadow : STD_ULOGIC;
signal V_E_CTRL_PC_shadow : PCTYPE;
signal V_E_CTRL_INST20_shadow : STD_LOGIC;
signal V_E_CTRL_WREG_shadow : STD_ULOGIC;
signal V_A_CTRL_WREG_shadow : STD_ULOGIC;
signal V_A_CTRL_shadow : PIPELINE_CTRL_TYPE;
signal V_A_CTRL_RD6DOWNTO0_shadow : std_logic_vector(6 downto 0);
signal V_X_DATA0_shadow : std_logic_vector(31 downto 0);
signal V_E_CTRL_INST19_shadow : STD_LOGIC;
signal ME_SIGNED_shadow : STD_ULOGIC;
signal V_W_WREG_shadow : STD_ULOGIC;
signal V_D_PC_shadow : PCTYPE;
signal VFPI_D_ANNUL_shadow : STD_ULOGIC;
signal DE_RADDR27DOWNTO0_shadow : STD_LOGIC_VECTOR(7 downto 0);
signal V_E_CTRL_CNT_shadow : OP_TYPE;
signal V_F_PC_shadow : PCTYPE;
signal V_X_DATA031_shadow : STD_LOGIC;
signal V_M_CTRL_PC31DOWNTO12_shadow : std_logic_vector(31 downto 12);
signal V_X_CTRL_RD7DOWNTO0_shadow : std_logic_vector(7 downto 0);
signal V_M_CTRL_TT_shadow : OP3_TYPE;
signal V_X_CTRL_shadow : PIPELINE_CTRL_TYPE;
signal V_A_CTRL_INST24_shadow : STD_LOGIC;
signal XC_TRAP_ADDRESS3DOWNTO2_shadow : std_logic_vector(3 downto 2);
signal V_X_NERROR_shadow : STD_ULOGIC;
signal V_F_PC31DOWNTO4_shadow : std_logic_vector(31 downto 4);
signal V_W_S_TT3DOWNTO0_shadow : STD_LOGIC_VECTOR(3 downto 0);
signal EX_JUMP_ADDRESS31DOWNTO4_shadow : std_logic_vector(31 downto 4);
signal EX_ADD_RES32DOWNTO332DOWNTO3_shadow : STD_LOGIC_VECTOR(32 downto 3);
signal V_F_BRANCH_shadow : STD_ULOGIC;
signal V_A_CTRL_WICC_shadow : STD_ULOGIC;
signal V_A_CTRL_LD_shadow : STD_ULOGIC;
signal V_A_CTRL_TT_shadow : OP3_TYPE;
signal V_M_CTRL_LD_shadow : STD_ULOGIC;
signal V_E_SHCNT_shadow : ASI_TYPE;
signal XC_TRAP_ADDRESS31DOWNTO12_shadow : std_logic_vector(31 downto 12);
signal V_A_CTRL_INST_shadow : WORD;
signal V_A_CTRL_RD7DOWNTO0_shadow : std_logic_vector(7 downto 0);
signal VIR_PWD_shadow : STD_ULOGIC;
signal XC_RESULT_shadow : WORD;
signal V_A_RFA1_shadow : RFATYPE;
signal V_E_JMPL_shadow : STD_ULOGIC;
signal V_E_CTRL_RD7DOWNTO0_shadow : std_logic_vector(7 downto 0);
signal ME_ICC_shadow : STD_LOGIC_VECTOR(3 downto 0);
signal DE_INST24_shadow : STD_LOGIC;
signal XC_TRAP_shadow : STD_ULOGIC;
signal VDSU_TBUFCNT_shadow : STD_LOGIC_VECTOR(6 downto 0);
signal XC_TRAP_ADDRESS_shadow : PCTYPE;

-- Intermediate value holding signal declarations
signal V_E_CTRL_WREG_shadow_intermed_2 : STD_ULOGIC;
signal V_M_CTRL_PC_shadow_intermed_2 : std_logic_vector(31 downto 2);
signal RIN_E_CTRL_TT3DOWNTO0_intermed_1 : std_logic_vector(3 downto 0);
signal V_D_PC3DOWNTO2_shadow_intermed_6 : std_logic_vector(3 downto 2);
signal RIN_M_CTRL_PC31DOWNTO12_intermed_5 : std_logic_vector(31 downto 12);
signal RIN_A_RFA1_intermed_1 : std_logic_vector(7 downto 0);
signal RIN_A_CTRL_PC31DOWNTO2_intermed_4 : std_logic_vector(31 downto 2);
signal R_E_CTRL_TT_intermed_1 : std_logic_vector(5 downto 0);
signal V_D_PC3DOWNTO2_shadow_intermed_2 : std_logic_vector(3 downto 2);
signal ICO_MEXC_intermed_4 : STD_ULOGIC;
signal V_F_PC31DOWNTO2_shadow_intermed_1 : std_logic_vector(31 downto 2);
signal RIN_X_DATA00_intermed_2 : STD_LOGIC;
signal R_A_CTRL_RD6DOWNTO0_intermed_1 : std_logic_vector(6 downto 0);
signal R_A_CTRL_INST24_intermed_1 : STD_LOGIC;
signal RIN_E_CTRL_INST19_intermed_1 : STD_LOGIC;
signal V_X_DATA00_shadow_intermed_3 : STD_LOGIC;
signal RIN_A_CTRL_INST19_intermed_2 : STD_LOGIC;
signal IRIN_ADDR31DOWNTO2_intermed_2 : std_logic_vector(31 downto 2);
signal V_E_CTRL_WREG_shadow_intermed_1 : STD_ULOGIC;
signal V_A_CTRL_PC31DOWNTO2_shadow_intermed_5 : std_logic_vector(31 downto 2);
signal V_M_CTRL_PC_shadow_intermed_3 : std_logic_vector(31 downto 2);
signal RIN_A_CTRL_WICC_intermed_3 : STD_ULOGIC;
signal V_A_CTRL_RETT_shadow_intermed_3 : STD_ULOGIC;
signal RPIN_PWD_intermed_1 : STD_ULOGIC;
signal RIN_A_CTRL_PC31DOWNTO12_intermed_7 : std_logic_vector(31 downto 12);
signal V_E_CTRL_TT_shadow_intermed_3 : std_logic_vector(5 downto 0);
signal DE_INST_shadow_intermed_2 : std_logic_vector(31 downto 0);
signal R_M_CTRL_PC31DOWNTO2_intermed_3 : std_logic_vector(31 downto 2);
signal DBGI_DADDR9DOWNTO2_intermed_1 : STD_LOGIC_VECTOR(9 downto 2);
signal R_D_PC31DOWNTO2_intermed_6 : std_logic_vector(31 downto 2);
signal RIN_A_CTRL_TT3DOWNTO0_intermed_5 : std_logic_vector(3 downto 0);
signal RIN_A_CTRL_TRAP_intermed_3 : STD_ULOGIC;
signal V_E_CTRL_CNT_shadow_intermed_2 : std_logic_vector(1 downto 0);
signal V_E_CTRL_PC31DOWNTO4_shadow_intermed_4 : std_logic_vector(31 downto 4);
signal RIN_D_STEP_intermed_1 : STD_ULOGIC;
signal V_M_CTRL_TT3DOWNTO0_shadow_intermed_4 : std_logic_vector(3 downto 0);
signal V_A_CTRL_PC_shadow_intermed_2 : std_logic_vector(31 downto 2);
signal RIN_D_PC31DOWNTO2_intermed_1 : std_logic_vector(31 downto 2);
signal V_E_CTRL_PC31DOWNTO4_shadow_intermed_5 : std_logic_vector(31 downto 4);
signal RIN_E_CTRL_INST20_intermed_1 : STD_LOGIC;
signal V_D_PC3DOWNTO2_shadow_intermed_7 : std_logic_vector(3 downto 2);
signal V_M_CTRL_PC31DOWNTO4_shadow_intermed_4 : std_logic_vector(31 downto 4);
signal V_M_CTRL_RD6DOWNTO0_shadow_intermed_2 : std_logic_vector(6 downto 0);
signal RIN_E_CTRL_PC3DOWNTO2_intermed_3 : std_logic_vector(3 downto 2);
signal RIN_M_Y31_intermed_1 : STD_LOGIC;
signal V_D_INST0_shadow_intermed_1 : std_logic_vector(31 downto 0);
signal RIN_E_YMSB_intermed_1 : STD_ULOGIC;
signal R_X_DATA031_intermed_2 : STD_LOGIC;
signal RIN_M_CTRL_WREG_intermed_2 : STD_ULOGIC;
signal V_X_CTRL_TT_shadow_intermed_1 : std_logic_vector(5 downto 0);
signal RIN_E_CTRL_PC_intermed_4 : std_logic_vector(31 downto 2);
signal V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2 : std_logic_vector(3 downto 0);
signal RIN_E_CTRL_PC31DOWNTO12_intermed_4 : std_logic_vector(31 downto 12);
signal V_A_CTRL_PC3DOWNTO2_shadow_intermed_3 : std_logic_vector(3 downto 2);
signal RIN_E_CTRL_PC31DOWNTO2_intermed_4 : std_logic_vector(31 downto 2);
signal R_A_CTRL_TT_intermed_1 : std_logic_vector(5 downto 0);
signal RIN_A_CTRL_WICC_intermed_2 : STD_ULOGIC;
signal V_E_CTRL_PC31DOWNTO2_shadow_intermed_6 : std_logic_vector(31 downto 2);
signal RIN_F_PC3DOWNTO2_intermed_1 : std_logic_vector(3 downto 2);
signal V_A_CTRL_PC31DOWNTO12_shadow_intermed_4 : std_logic_vector(31 downto 12);
signal EX_ADD_RES32DOWNTO332DOWNTO5_shadow_intermed_1 : STD_LOGIC_VECTOR(32 downto 5);
signal V_X_DATA04DOWNTO0_shadow_intermed_1 : std_logic_vector(4 downto 0);
signal R_A_CTRL_INST20_intermed_2 : STD_LOGIC;
signal V_A_CTRL_PC31DOWNTO12_shadow_intermed_6 : std_logic_vector(31 downto 12);
signal R_A_CTRL_RETT_intermed_2 : STD_ULOGIC;
signal RIN_M_DCI_LOCK_intermed_1 : STD_ULOGIC;
signal RIN_D_PC31DOWNTO12_intermed_6 : std_logic_vector(31 downto 12);
signal RIN_E_CTRL_TT_intermed_3 : std_logic_vector(5 downto 0);
signal R_E_CTRL_RD7DOWNTO0_intermed_2 : std_logic_vector(7 downto 0);
signal RIN_A_ET_intermed_1 : STD_ULOGIC;
signal RIN_X_CTRL_RD6DOWNTO0_intermed_1 : std_logic_vector(6 downto 0);
signal RIN_M_CTRL_PC31DOWNTO12_intermed_2 : std_logic_vector(31 downto 12);
signal DBGI_STEP_intermed_1 : STD_ULOGIC;
signal V_A_CTRL_RETT_shadow_intermed_2 : STD_ULOGIC;
signal R_X_CTRL_PC3DOWNTO2_intermed_1 : std_logic_vector(3 downto 2);
signal R_A_CTRL_PC31DOWNTO4_intermed_4 : std_logic_vector(31 downto 4);
signal V_M_CTRL_PV_shadow_intermed_1 : STD_ULOGIC;
signal RIN_M_CTRL_PC31DOWNTO2_intermed_5 : std_logic_vector(31 downto 2);
signal V_M_CTRL_PC31DOWNTO12_shadow_intermed_5 : std_logic_vector(31 downto 12);
signal V_X_LADDR_shadow_intermed_1 : std_logic_vector(1 downto 0);
signal V_D_ANNUL_shadow_intermed_2 : STD_ULOGIC;
signal V_A_CTRL_RD6DOWNTO0_shadow_intermed_1 : std_logic_vector(6 downto 0);
signal RIN_W_WA_intermed_1 : std_logic_vector(7 downto 0);
signal V_D_PC_shadow_intermed_4 : std_logic_vector(31 downto 2);
signal V_X_CTRL_PC31DOWNTO2_shadow_intermed_1 : std_logic_vector(31 downto 2);
signal RIN_X_CTRL_PC31DOWNTO4_intermed_2 : std_logic_vector(31 downto 4);
signal V_E_CTRL_WICC_shadow_intermed_1 : STD_ULOGIC;
signal VDSU_CRDY2_shadow_intermed_2 : STD_LOGIC;
signal V_M_RESULT1DOWNTO0_shadow_intermed_3 : std_logic_vector(1 downto 0);
signal RIN_D_INST0_intermed_1 : std_logic_vector(31 downto 0);
signal V_X_DATA03_shadow_intermed_2 : STD_LOGIC;
signal RIN_X_DCI_intermed_1 : DC_IN_TYPE;
signal DSUIN_TT_intermed_1 : STD_LOGIC_VECTOR(7 downto 0);
signal V_D_CNT_shadow_intermed_4 : std_logic_vector(1 downto 0);
signal RIN_D_CNT_intermed_4 : std_logic_vector(1 downto 0);
signal ICO_MEXC_intermed_1 : STD_ULOGIC;
signal R_X_ANNUL_ALL_intermed_2 : STD_ULOGIC;
signal R_X_CTRL_TT3DOWNTO0_intermed_2 : std_logic_vector(3 downto 0);
signal R_D_PC3DOWNTO2_intermed_3 : std_logic_vector(3 downto 2);
signal RIN_D_CNT_intermed_2 : std_logic_vector(1 downto 0);
signal V_M_DCI_SIZE_shadow_intermed_2 : std_logic_vector(1 downto 0);
signal R_A_CTRL_ANNUL_intermed_2 : STD_ULOGIC;
signal V_W_S_S_shadow_intermed_1 : STD_ULOGIC;
signal RIN_M_CTRL_TT_intermed_2 : std_logic_vector(5 downto 0);
signal EX_ADD_RES32DOWNTO330DOWNTO11_shadow_intermed_1 : STD_LOGIC_VECTOR(30 downto 11);
signal V_A_CTRL_RETT_shadow_intermed_1 : STD_ULOGIC;
signal R_X_DATA04DOWNTO0_intermed_1 : std_logic_vector(4 downto 0);
signal V_E_CTRL_TT3DOWNTO0_shadow_intermed_1 : std_logic_vector(3 downto 0);
signal V_D_PC31DOWNTO4_shadow_intermed_6 : std_logic_vector(31 downto 4);
signal V_X_CTRL_RD6DOWNTO0_shadow_intermed_1 : std_logic_vector(6 downto 0);
signal RIN_W_S_ET_intermed_1 : STD_ULOGIC;
signal R_E_CTRL_TRAP_intermed_1 : STD_ULOGIC;
signal V_A_CTRL_PC_shadow_intermed_3 : std_logic_vector(31 downto 2);
signal R_M_CTRL_PC31DOWNTO4_intermed_2 : std_logic_vector(31 downto 4);
signal VIR_ADDR31DOWNTO4_shadow_intermed_2 : std_logic_vector(31 downto 4);
signal V_E_CTRL_RD6DOWNTO0_shadow_intermed_3 : std_logic_vector(6 downto 0);
signal R_D_CWP_intermed_1 : std_logic_vector(2 downto 0);
signal RIN_A_CTRL_TT3DOWNTO0_intermed_2 : std_logic_vector(3 downto 0);
signal RIN_X_CTRL_PC3DOWNTO2_intermed_3 : std_logic_vector(3 downto 2);
signal RIN_D_PC31DOWNTO2_intermed_8 : std_logic_vector(31 downto 2);
signal RIN_A_CTRL_ANNUL_intermed_1 : STD_ULOGIC;
signal V_X_CTRL_PC3DOWNTO2_shadow_intermed_1 : std_logic_vector(3 downto 2);
signal RIN_M_CTRL_PC31DOWNTO12_intermed_3 : std_logic_vector(31 downto 12);
signal R_M_DCI_SIGNED_intermed_1 : STD_ULOGIC;
signal RIN_X_DCI_SIGNED_intermed_1 : STD_ULOGIC;
signal V_D_PC31DOWNTO2_shadow_intermed_4 : std_logic_vector(31 downto 2);
signal DCO_DATA00_intermed_2 : STD_LOGIC;
signal V_M_CTRL_RD7DOWNTO0_shadow_intermed_2 : std_logic_vector(7 downto 0);
signal V_E_SU_shadow_intermed_1 : STD_ULOGIC;
signal R_A_CTRL_INST20_intermed_1 : STD_LOGIC;
signal R_D_PC31DOWNTO12_intermed_7 : std_logic_vector(31 downto 12);
signal XC_TRAP_ADDRESS_shadow_intermed_1 : std_logic_vector(31 downto 2);
signal RIN_X_CTRL_PC31DOWNTO2_intermed_3 : std_logic_vector(31 downto 2);
signal R_E_CTRL_RETT_intermed_1 : STD_ULOGIC;
signal V_X_DCI_SIZE_shadow_intermed_1 : std_logic_vector(1 downto 0);
signal RIN_D_CNT_intermed_3 : std_logic_vector(1 downto 0);
signal RIN_A_CTRL_ANNUL_intermed_4 : STD_ULOGIC;
signal R_E_CTRL_TT3DOWNTO0_intermed_1 : std_logic_vector(3 downto 0);
signal R_D_PC3DOWNTO2_intermed_2 : std_logic_vector(3 downto 2);
signal V_X_CTRL_TT3DOWNTO0_shadow_intermed_3 : std_logic_vector(3 downto 0);
signal V_A_CTRL_RD6DOWNTO0_shadow_intermed_3 : std_logic_vector(6 downto 0);
signal R_M_CTRL_PC31DOWNTO2_intermed_4 : std_logic_vector(31 downto 2);
signal RIN_A_CTRL_PC31DOWNTO12_intermed_3 : std_logic_vector(31 downto 12);
signal R_A_CTRL_PC31DOWNTO12_intermed_5 : std_logic_vector(31 downto 12);
signal R_A_CTRL_PC_intermed_2 : std_logic_vector(31 downto 2);
signal V_X_MEXC_shadow_intermed_1 : STD_ULOGIC;
signal V_M_CTRL_RD7DOWNTO0_shadow_intermed_1 : std_logic_vector(7 downto 0);
signal IR_ADDR31DOWNTO4_intermed_1 : std_logic_vector(31 downto 4);
signal V_A_CTRL_PC_shadow_intermed_4 : std_logic_vector(31 downto 2);
signal VIR_ADDR31DOWNTO4_shadow_intermed_1 : std_logic_vector(31 downto 4);
signal RIN_M_CTRL_PC3DOWNTO2_intermed_1 : std_logic_vector(3 downto 2);
signal RIN_E_CTRL_WREG_intermed_1 : STD_ULOGIC;
signal RIN_D_PC31DOWNTO12_intermed_1 : std_logic_vector(31 downto 12);
signal V_E_CTRL_TT3DOWNTO0_shadow_intermed_2 : std_logic_vector(3 downto 0);
signal RIN_D_INST1_intermed_1 : std_logic_vector(31 downto 0);
signal RIN_D_PC31DOWNTO12_intermed_3 : std_logic_vector(31 downto 12);
signal V_A_CTRL_TT_shadow_intermed_3 : std_logic_vector(5 downto 0);
signal RIN_A_CTRL_INST24_intermed_2 : STD_LOGIC;
signal V_X_DATA1_shadow_intermed_2 : std_logic_vector(31 downto 0);
signal ICO_MEXC_intermed_3 : STD_ULOGIC;
signal R_D_PC3DOWNTO2_intermed_4 : std_logic_vector(3 downto 2);
signal R_M_CTRL_INST_intermed_1 : std_logic_vector(31 downto 0);
signal V_A_CWP_shadow_intermed_1 : std_logic_vector(2 downto 0);
signal V_A_CTRL_WICC_shadow_intermed_3 : STD_ULOGIC;
signal V_D_PC_shadow_intermed_6 : std_logic_vector(31 downto 2);
signal RIN_X_ANNUL_ALL_intermed_5 : STD_ULOGIC;
signal RIN_E_CTRL_INST20_intermed_2 : STD_LOGIC;
signal R_X_DATA0_intermed_2 : std_logic_vector(31 downto 0);
signal RIN_D_PC_intermed_4 : std_logic_vector(31 downto 2);
signal R_E_CTRL_PV_intermed_1 : STD_ULOGIC;
signal R_E_CTRL_TT3DOWNTO0_intermed_2 : std_logic_vector(3 downto 0);
signal R_D_PC_intermed_1 : std_logic_vector(31 downto 2);
signal R_A_CTRL_PC_intermed_3 : std_logic_vector(31 downto 2);
signal EX_JUMP_ADDRESS31DOWNTO12_shadow_intermed_1 : std_logic_vector(31 downto 12);
signal R_X_CTRL_TT3DOWNTO0_intermed_1 : std_logic_vector(3 downto 0);
signal V_M_DCI_SIGNED_shadow_intermed_1 : STD_ULOGIC;
signal RIN_X_CTRL_TT3DOWNTO0_intermed_1 : std_logic_vector(3 downto 0);
signal V_X_ANNUL_ALL_shadow_intermed_2 : STD_ULOGIC;
signal V_D_PC31DOWNTO4_shadow_intermed_7 : std_logic_vector(31 downto 4);
signal RIN_E_OP13_intermed_1 : STD_LOGIC;
signal RIN_A_CWP_intermed_1 : std_logic_vector(2 downto 0);
signal RIN_E_CTRL_WICC_intermed_1 : STD_ULOGIC;
signal VP_ERROR_shadow_intermed_2 : STD_ULOGIC;
signal RIN_E_OP2_intermed_1 : std_logic_vector(31 downto 0);
signal RIN_A_CTRL_TT3DOWNTO0_intermed_4 : std_logic_vector(3 downto 0);
signal RIN_A_CTRL_RD7DOWNTO0_intermed_2 : std_logic_vector(7 downto 0);
signal RIN_E_CTRL_intermed_2 : PIPELINE_CTRL_TYPE;
signal R_M_CTRL_PC_intermed_1 : std_logic_vector(31 downto 2);
signal RIN_E_CTRL_PC31DOWNTO2_intermed_5 : std_logic_vector(31 downto 2);
signal R_M_Y31_intermed_2 : STD_LOGIC;
signal V_M_CTRL_PC3DOWNTO2_shadow_intermed_4 : std_logic_vector(3 downto 2);
signal V_M_CTRL_RETT_shadow_intermed_1 : STD_ULOGIC;
signal V_X_CTRL_PC31DOWNTO4_shadow_intermed_3 : std_logic_vector(31 downto 4);
signal XC_VECTT3DOWNTO0_shadow_intermed_2 : STD_LOGIC_VECTOR(3 downto 0);
signal RIN_M_CTRL_PC31DOWNTO12_intermed_1 : std_logic_vector(31 downto 12);
signal RIN_M_RESULT1DOWNTO0_intermed_2 : std_logic_vector(1 downto 0);
signal V_X_ANNUL_ALL_shadow_intermed_4 : STD_ULOGIC;
signal RIN_W_S_TBA_intermed_1 : STD_LOGIC_VECTOR(19 downto 0);
signal V_D_INST1_shadow_intermed_1 : std_logic_vector(31 downto 0);
signal RIN_X_DATA031_intermed_1 : STD_LOGIC;
signal XC_TRAP_ADDRESS31DOWNTO12_shadow_intermed_1 : std_logic_vector(31 downto 12);
signal RIN_D_PC3DOWNTO2_intermed_4 : std_logic_vector(3 downto 2);
signal RIN_X_CTRL_PC31DOWNTO4_intermed_3 : std_logic_vector(31 downto 4);
signal V_E_CTRL_PC31DOWNTO4_shadow_intermed_2 : std_logic_vector(31 downto 4);
signal V_M_CTRL_PC3DOWNTO2_shadow_intermed_3 : std_logic_vector(3 downto 2);
signal V_M_CTRL_PC31DOWNTO12_shadow_intermed_2 : std_logic_vector(31 downto 12);
signal RIN_E_CTRL_PV_intermed_1 : STD_ULOGIC;
signal EX_ADD_RES32DOWNTO332DOWNTO13_shadow_intermed_1 : STD_LOGIC_VECTOR(32 downto 13);
signal R_E_CTRL_WREG_intermed_2 : STD_ULOGIC;
signal R_X_DATA031_intermed_1 : STD_LOGIC;
signal R_D_INST0_intermed_2 : std_logic_vector(31 downto 0);
signal RIN_E_SARI_intermed_1 : STD_ULOGIC;
signal R_M_Y31_intermed_1 : STD_LOGIC;
signal IR_ADDR3DOWNTO2_intermed_1 : std_logic_vector(3 downto 2);
signal DE_INST24_shadow_intermed_2 : STD_LOGIC;
signal V_W_S_S_shadow_intermed_2 : STD_ULOGIC;
signal DE_INST20_shadow_intermed_3 : STD_LOGIC;
signal R_E_CTRL_TT3DOWNTO0_intermed_4 : std_logic_vector(3 downto 0);
signal RIN_A_CTRL_TT_intermed_2 : std_logic_vector(5 downto 0);
signal V_A_CTRL_PV_shadow_intermed_2 : STD_ULOGIC;
signal V_E_CTRL_TT_shadow_intermed_1 : std_logic_vector(5 downto 0);
signal V_D_PC31DOWNTO2_shadow_intermed_5 : std_logic_vector(31 downto 2);
signal V_X_DATA04DOWNTO0_shadow_intermed_2 : std_logic_vector(4 downto 0);
signal R_X_CTRL_PC31DOWNTO4_intermed_2 : std_logic_vector(31 downto 4);
signal RIN_M_CTRL_INST_intermed_1 : std_logic_vector(31 downto 0);
signal RIN_A_CTRL_RD6DOWNTO0_intermed_2 : std_logic_vector(6 downto 0);
signal DCO_DATA04DOWNTO0_intermed_2 : std_logic_vector(4 downto 0);
signal EX_JUMP_ADDRESS31DOWNTO12_shadow_intermed_2 : std_logic_vector(31 downto 12);
signal V_X_DATA0_shadow_intermed_2 : std_logic_vector(31 downto 0);
signal R_A_CTRL_WREG_intermed_3 : STD_ULOGIC;
signal RIN_X_CTRL_PC31DOWNTO12_intermed_2 : std_logic_vector(31 downto 12);
signal R_D_CNT_intermed_3 : std_logic_vector(1 downto 0);
signal V_E_OP131_shadow_intermed_1 : STD_LOGIC;
signal R_D_PC31DOWNTO12_intermed_6 : std_logic_vector(31 downto 12);
signal RIN_X_CTRL_WICC_intermed_1 : STD_ULOGIC;
signal V_D_PC31DOWNTO12_shadow_intermed_1 : std_logic_vector(31 downto 12);
signal RIN_E_CTRL_TRAP_intermed_3 : STD_ULOGIC;
signal R_X_RESULT6DOWNTO0_intermed_1 : std_logic_vector(6 downto 0);
signal R_E_CTRL_INST19_intermed_2 : STD_LOGIC;
signal RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2 : std_logic_vector(3 downto 0);
signal R_M_CTRL_RD7DOWNTO0_intermed_1 : std_logic_vector(7 downto 0);
signal RIN_E_CTRL_PC31DOWNTO12_intermed_6 : std_logic_vector(31 downto 12);
signal RIN_A_CTRL_PC31DOWNTO4_intermed_3 : std_logic_vector(31 downto 4);
signal V_A_CTRL_INST19_shadow_intermed_3 : STD_LOGIC;
signal V_D_PC31DOWNTO12_shadow_intermed_5 : std_logic_vector(31 downto 12);
signal V_A_CTRL_INST19_shadow_intermed_2 : STD_LOGIC;
signal V_X_CTRL_WREG_shadow_intermed_1 : STD_ULOGIC;
signal V_A_CTRL_TRAP_shadow_intermed_2 : STD_ULOGIC;
signal RIN_E_CTRL_PC3DOWNTO2_intermed_1 : std_logic_vector(3 downto 2);
signal RIN_M_CTRL_PC3DOWNTO2_intermed_3 : std_logic_vector(3 downto 2);
signal V_A_RFE2_shadow_intermed_1 : STD_ULOGIC;
signal V_M_Y_shadow_intermed_1 : std_logic_vector(31 downto 0);
signal RIN_A_CTRL_LD_intermed_1 : STD_ULOGIC;
signal V_E_CTRL_PC_shadow_intermed_3 : std_logic_vector(31 downto 2);
signal RIN_D_INST1_intermed_2 : std_logic_vector(31 downto 0);
signal R_E_CTRL_PC31DOWNTO12_intermed_1 : std_logic_vector(31 downto 12);
signal RIN_X_CTRL_PC31DOWNTO12_intermed_3 : std_logic_vector(31 downto 12);
signal R_E_CTRL_TRAP_intermed_2 : STD_ULOGIC;
signal DE_INST24_shadow_intermed_1 : STD_LOGIC;
signal V_E_CTRL_PC_shadow_intermed_2 : std_logic_vector(31 downto 2);
signal V_A_CTRL_TT_shadow_intermed_1 : std_logic_vector(5 downto 0);
signal V_D_MEXC_shadow_intermed_4 : STD_ULOGIC;
signal V_D_PC31DOWNTO12_shadow_intermed_6 : std_logic_vector(31 downto 12);
signal V_A_CTRL_PC31DOWNTO12_shadow_intermed_3 : std_logic_vector(31 downto 12);
signal R_X_CTRL_PC31DOWNTO12_intermed_3 : std_logic_vector(31 downto 12);
signal V_M_CTRL_PV_shadow_intermed_2 : STD_ULOGIC;
signal RIN_A_CTRL_PC31DOWNTO2_intermed_2 : std_logic_vector(31 downto 2);
signal EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_2 : std_logic_vector(31 downto 2);
signal RIN_E_CTRL_PC31DOWNTO4_intermed_1 : std_logic_vector(31 downto 4);
signal RIN_E_CTRL_PC31DOWNTO12_intermed_2 : std_logic_vector(31 downto 12);
signal RIN_M_CTRL_TRAP_intermed_1 : STD_ULOGIC;
signal R_E_CTRL_PC31DOWNTO2_intermed_2 : std_logic_vector(31 downto 2);
signal R_E_CTRL_LD_intermed_1 : STD_ULOGIC;
signal R_M_CTRL_PC31DOWNTO2_intermed_1 : std_logic_vector(31 downto 2);
signal RIN_A_CTRL_PC31DOWNTO2_intermed_5 : std_logic_vector(31 downto 2);
signal V_W_S_CWP_shadow_intermed_1 : std_logic_vector(2 downto 0);
signal R_M_CTRL_PC3DOWNTO2_intermed_1 : std_logic_vector(3 downto 2);
signal V_E_CTRL_PC31DOWNTO12_shadow_intermed_4 : std_logic_vector(31 downto 12);
signal R_X_CTRL_PC31DOWNTO4_intermed_1 : std_logic_vector(31 downto 4);
signal V_M_CTRL_PC_shadow_intermed_1 : std_logic_vector(31 downto 2);
signal IR_ADDR31DOWNTO2_intermed_2 : std_logic_vector(31 downto 2);
signal V_E_CTRL_TT3DOWNTO0_shadow_intermed_4 : std_logic_vector(3 downto 0);
signal V_E_CTRL_PC3DOWNTO2_shadow_intermed_3 : std_logic_vector(3 downto 2);
signal RIN_X_CTRL_PC31DOWNTO4_intermed_1 : std_logic_vector(31 downto 4);
signal R_E_CTRL_PC31DOWNTO12_intermed_2 : std_logic_vector(31 downto 12);
signal RIN_M_CTRL_RETT_intermed_1 : STD_ULOGIC;
signal V_M_DCI_LOCK_shadow_intermed_1 : STD_ULOGIC;
signal V_X_RESULT6DOWNTO0_shadow_intermed_1 : std_logic_vector(6 downto 0);
signal RIN_X_DATA04DOWNTO0_intermed_3 : std_logic_vector(4 downto 0);
signal V_X_NERROR_shadow_intermed_1 : STD_ULOGIC;
signal V_A_RFE1_shadow_intermed_1 : STD_ULOGIC;
signal V_D_PC3DOWNTO2_shadow_intermed_1 : std_logic_vector(3 downto 2);
signal V_E_CTRL_LD_shadow_intermed_1 : STD_ULOGIC;
signal ICO_DATA0_intermed_1 : std_logic_vector(31 downto 0);
signal VIR_ADDR_shadow_intermed_1 : std_logic_vector(31 downto 2);
signal R_M_CTRL_PC31DOWNTO12_intermed_2 : std_logic_vector(31 downto 12);
signal V_E_CTRL_PV_shadow_intermed_2 : STD_ULOGIC;
signal RIN_E_CTRL_PC31DOWNTO4_intermed_4 : std_logic_vector(31 downto 4);
signal R_A_CTRL_PC3DOWNTO2_intermed_3 : std_logic_vector(3 downto 2);
signal R_E_CTRL_INST19_intermed_1 : STD_LOGIC;
signal RIN_E_CTRL_TT3DOWNTO0_intermed_4 : std_logic_vector(3 downto 0);
signal R_M_CTRL_PC31DOWNTO4_intermed_3 : std_logic_vector(31 downto 4);
signal V_A_CTRL_PC31DOWNTO4_shadow_intermed_4 : std_logic_vector(31 downto 4);
signal RIN_W_S_DWT_intermed_1 : STD_ULOGIC;
signal V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 : std_logic_vector(31 downto 2);
signal R_D_PC31DOWNTO12_intermed_4 : std_logic_vector(31 downto 12);
signal RIN_X_NERROR_intermed_1 : STD_ULOGIC;
signal R_M_CTRL_PC3DOWNTO2_intermed_2 : std_logic_vector(3 downto 2);
signal ICO_MEXC_intermed_5 : STD_ULOGIC;
signal R_A_CTRL_RD7DOWNTO0_intermed_2 : std_logic_vector(7 downto 0);
signal V_A_CTRL_PC31DOWNTO4_shadow_intermed_1 : std_logic_vector(31 downto 4);
signal IRIN_ADDR31DOWNTO2_intermed_1 : std_logic_vector(31 downto 2);
signal VIR_ADDR31DOWNTO12_shadow_intermed_3 : std_logic_vector(31 downto 12);
signal XC_TRAP_ADDRESS3DOWNTO2_shadow_intermed_1 : std_logic_vector(3 downto 2);
signal R_A_CTRL_INST_intermed_1 : std_logic_vector(31 downto 0);
signal R_E_CTRL_PC31DOWNTO2_intermed_3 : std_logic_vector(31 downto 2);
signal RIN_X_CTRL_TT3DOWNTO0_intermed_3 : std_logic_vector(3 downto 0);
signal RIN_M_CTRL_PC3DOWNTO2_intermed_2 : std_logic_vector(3 downto 2);
signal V_M_CTRL_PC31DOWNTO2_shadow_intermed_4 : std_logic_vector(31 downto 2);
signal RIN_A_CTRL_RETT_intermed_2 : STD_ULOGIC;
signal V_X_DATA00_shadow_intermed_1 : STD_LOGIC;
signal RIN_M_CTRL_RD6DOWNTO0_intermed_2 : std_logic_vector(6 downto 0);
signal RIN_E_CTRL_TT3DOWNTO0_intermed_2 : std_logic_vector(3 downto 0);
signal V_M_CTRL_INST_shadow_intermed_1 : std_logic_vector(31 downto 0);
signal RIN_A_CTRL_TT3DOWNTO0_intermed_3 : std_logic_vector(3 downto 0);
signal EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_1 : STD_LOGIC_VECTOR(32 downto 3);
signal R_A_CTRL_TT3DOWNTO0_intermed_1 : std_logic_vector(3 downto 0);
signal V_X_DEBUG_shadow_intermed_1 : STD_ULOGIC;
signal V_E_CTRL_PC_shadow_intermed_4 : std_logic_vector(31 downto 2);
signal V_M_CTRL_TT_shadow_intermed_1 : std_logic_vector(5 downto 0);
signal RIN_A_CTRL_PV_intermed_4 : STD_ULOGIC;
signal R_E_MAC_intermed_1 : STD_ULOGIC;
signal V_E_CTRL_PC3DOWNTO2_shadow_intermed_1 : std_logic_vector(3 downto 2);
signal R_M_RESULT1DOWNTO0_intermed_1 : std_logic_vector(1 downto 0);
signal IR_ADDR31DOWNTO2_intermed_1 : std_logic_vector(31 downto 2);
signal RIN_A_CTRL_WREG_intermed_2 : STD_ULOGIC;
signal V_D_MEXC_shadow_intermed_1 : STD_ULOGIC;
signal XC_TRAP_ADDRESS31DOWNTO12_shadow_intermed_2 : std_logic_vector(31 downto 12);
signal R_A_CTRL_LD_intermed_2 : STD_ULOGIC;
signal R_A_CTRL_intermed_2 : PIPELINE_CTRL_TYPE;
signal V_M_CTRL_TRAP_shadow_intermed_2 : STD_ULOGIC;
signal V_A_JMPL_shadow_intermed_1 : STD_ULOGIC;
signal V_E_CTRL_RETT_shadow_intermed_2 : STD_ULOGIC;
signal RIN_M_CTRL_LD_intermed_1 : STD_ULOGIC;
signal V_X_DATA04DOWNTO0_shadow_intermed_3 : std_logic_vector(4 downto 0);
signal RIN_W_S_TT_intermed_1 : STD_LOGIC_VECTOR(7 downto 0);
signal V_A_CTRL_PC_shadow_intermed_5 : std_logic_vector(31 downto 2);
signal V_X_CTRL_PC31DOWNTO12_shadow_intermed_1 : std_logic_vector(31 downto 12);
signal DCO_DATA031_intermed_1 : STD_LOGIC;
signal RIN_A_CTRL_CNT_intermed_1 : std_logic_vector(1 downto 0);
signal R_X_ANNUL_ALL_intermed_3 : STD_ULOGIC;
signal V_X_DATA031_shadow_intermed_3 : STD_LOGIC;
signal DCO_DATA1_intermed_1 : std_logic_vector(31 downto 0);
signal V_E_CTRL_RETT_shadow_intermed_1 : STD_ULOGIC;
signal RIN_E_CTRL_CNT_intermed_1 : std_logic_vector(1 downto 0);
signal V_X_DATA0_shadow_intermed_1 : std_logic_vector(31 downto 0);
signal V_A_CTRL_LD_shadow_intermed_2 : STD_ULOGIC;
signal V_A_CTRL_TT3DOWNTO0_shadow_intermed_6 : std_logic_vector(3 downto 0);
signal R_E_CTRL_PC31DOWNTO4_intermed_3 : std_logic_vector(31 downto 4);
signal RPIN_ERROR_intermed_1 : STD_ULOGIC;
signal V_X_CTRL_PC31DOWNTO2_shadow_intermed_3 : std_logic_vector(31 downto 2);
signal R_W_S_S_intermed_1 : STD_ULOGIC;
signal R_A_CTRL_WICC_intermed_1 : STD_ULOGIC;
signal RIN_A_CTRL_PC31DOWNTO4_intermed_5 : std_logic_vector(31 downto 4);
signal RIN_D_PC31DOWNTO4_intermed_1 : std_logic_vector(31 downto 4);
signal EX_JUMP_ADDRESS31DOWNTO4_shadow_intermed_1 : std_logic_vector(31 downto 4);
signal RIN_D_PC_intermed_5 : std_logic_vector(31 downto 2);
signal V_A_RFA1_shadow_intermed_1 : std_logic_vector(7 downto 0);
signal R_X_CTRL_PC31DOWNTO2_intermed_1 : std_logic_vector(31 downto 2);
signal R_D_PC_intermed_2 : std_logic_vector(31 downto 2);
signal V_A_CTRL_PC3DOWNTO2_shadow_intermed_5 : std_logic_vector(3 downto 2);
signal RIN_E_SU_intermed_1 : STD_ULOGIC;
signal V_E_CTRL_INST_shadow_intermed_1 : std_logic_vector(31 downto 0);
signal RIN_M_CTRL_PC_intermed_1 : std_logic_vector(31 downto 2);
signal R_X_ANNUL_ALL_intermed_4 : STD_ULOGIC;
signal RIN_A_CTRL_INST_intermed_3 : std_logic_vector(31 downto 0);
signal V_A_CTRL_shadow_intermed_3 : PIPELINE_CTRL_TYPE;
signal R_D_MEXC_intermed_1 : STD_ULOGIC;
signal RIN_X_CTRL_RETT_intermed_1 : STD_ULOGIC;
signal R_X_RESULT6DOWNTO03DOWNTO0_intermed_1 : std_logic_vector(3 downto 0);
signal R_A_CTRL_WICC_intermed_2 : STD_ULOGIC;
signal VDSU_CRDY2_shadow_intermed_1 : STD_LOGIC;
signal V_A_DIVSTART_shadow_intermed_1 : STD_ULOGIC;
signal R_A_CTRL_PC31DOWNTO2_intermed_6 : std_logic_vector(31 downto 2);
signal RIN_A_CTRL_TRAP_intermed_4 : STD_ULOGIC;
signal RIN_W_S_PS_intermed_1 : STD_ULOGIC;
signal R_D_MEXC_intermed_3 : STD_ULOGIC;
signal RIN_A_RFA2_intermed_1 : std_logic_vector(7 downto 0);
signal R_X_DATA1_intermed_1 : std_logic_vector(31 downto 0);
signal V_A_CTRL_PV_shadow_intermed_1 : STD_ULOGIC;
signal R_A_CTRL_PC31DOWNTO4_intermed_1 : std_logic_vector(31 downto 4);
signal V_X_CTRL_PC31DOWNTO4_shadow_intermed_2 : std_logic_vector(31 downto 4);
signal RIN_W_S_SVT_intermed_1 : STD_ULOGIC;
signal RIN_E_CTRL_RD6DOWNTO0_intermed_1 : std_logic_vector(6 downto 0);
signal R_D_PC31DOWNTO12_intermed_5 : std_logic_vector(31 downto 12);
signal RIN_A_CTRL_INST19_intermed_1 : STD_LOGIC;
signal RIN_M_CTRL_PV_intermed_1 : STD_ULOGIC;
signal RIN_A_CTRL_RD6DOWNTO0_intermed_4 : std_logic_vector(6 downto 0);
signal RIN_E_OP23_intermed_1 : STD_LOGIC;
signal RIN_E_CTRL_WICC_intermed_2 : STD_ULOGIC;
signal R_D_PC31DOWNTO4_intermed_5 : std_logic_vector(31 downto 4);
signal V_D_MEXC_shadow_intermed_2 : STD_ULOGIC;
signal RIN_D_PC31DOWNTO4_intermed_7 : std_logic_vector(31 downto 4);
signal R_A_CTRL_TRAP_intermed_3 : STD_ULOGIC;
signal V_E_CTRL_INST19_shadow_intermed_2 : STD_LOGIC;
signal RIN_E_CTRL_PC31DOWNTO12_intermed_5 : std_logic_vector(31 downto 12);
signal RIN_D_PC31DOWNTO12_intermed_8 : std_logic_vector(31 downto 12);
signal VP_PWD_shadow_intermed_1 : STD_ULOGIC;
signal RIN_M_CTRL_RD7DOWNTO0_intermed_1 : std_logic_vector(7 downto 0);
signal V_A_CTRL_PC31DOWNTO4_shadow_intermed_2 : std_logic_vector(31 downto 4);
signal RIN_F_PC31DOWNTO2_intermed_2 : std_logic_vector(31 downto 2);
signal RIN_M_NALIGN_intermed_1 : STD_ULOGIC;
signal RP_ERROR_intermed_1 : STD_ULOGIC;
signal RIN_X_CTRL_PC3DOWNTO2_intermed_2 : std_logic_vector(3 downto 2);
signal V_W_S_TBA_shadow_intermed_1 : STD_LOGIC_VECTOR(19 downto 0);
signal R_F_PC31DOWNTO12_intermed_2 : std_logic_vector(31 downto 12);
signal RIN_E_JMPL_intermed_1 : STD_ULOGIC;
signal RIN_A_CTRL_TRAP_intermed_1 : STD_ULOGIC;
signal V_A_SU_shadow_intermed_1 : STD_ULOGIC;
signal RIN_A_RFE2_intermed_1 : STD_ULOGIC;
signal RIN_D_PC_intermed_2 : std_logic_vector(31 downto 2);
signal RIN_A_CTRL_CNT_intermed_3 : std_logic_vector(1 downto 0);
signal V_M_CTRL_PC31DOWNTO12_shadow_intermed_3 : std_logic_vector(31 downto 12);
signal V_M_CTRL_PC3DOWNTO2_shadow_intermed_2 : std_logic_vector(3 downto 2);
signal VIR_ADDR31DOWNTO12_shadow_intermed_1 : std_logic_vector(31 downto 12);
signal RIN_E_CTRL_LD_intermed_2 : STD_ULOGIC;
signal V_E_CTRL_PC31DOWNTO12_shadow_intermed_2 : std_logic_vector(31 downto 12);
signal R_E_CTRL_PC31DOWNTO12_intermed_4 : std_logic_vector(31 downto 12);
signal V_X_CTRL_PC3DOWNTO2_shadow_intermed_2 : std_logic_vector(3 downto 2);
signal V_A_CTRL_INST24_shadow_intermed_2 : STD_LOGIC;
signal V_M_CTRL_TRAP_shadow_intermed_1 : STD_ULOGIC;
signal V_E_CTRL_PC31DOWNTO4_shadow_intermed_3 : std_logic_vector(31 downto 4);
signal V_A_CTRL_PC3DOWNTO2_shadow_intermed_4 : std_logic_vector(3 downto 2);
signal R_A_CTRL_PC31DOWNTO2_intermed_5 : std_logic_vector(31 downto 2);
signal R_X_DATA0_intermed_1 : std_logic_vector(31 downto 0);
signal V_E_CTRL_TT_shadow_intermed_2 : std_logic_vector(5 downto 0);
signal V_E_MAC_shadow_intermed_2 : STD_ULOGIC;
signal RIN_E_CTRL_INST19_intermed_2 : STD_LOGIC;
signal RIN_D_PC31DOWNTO2_intermed_3 : std_logic_vector(31 downto 2);
signal IRIN_ADDR_intermed_1 : std_logic_vector(31 downto 2);
signal RIN_X_ANNUL_ALL_intermed_3 : STD_ULOGIC;
signal RIN_E_CTRL_INST_intermed_2 : std_logic_vector(31 downto 0);
signal V_X_CTRL_PC_shadow_intermed_2 : std_logic_vector(31 downto 2);
signal R_M_CTRL_TRAP_intermed_1 : STD_ULOGIC;
signal V_D_CWP_shadow_intermed_2 : std_logic_vector(2 downto 0);
signal V_A_CTRL_PC31DOWNTO12_shadow_intermed_2 : std_logic_vector(31 downto 12);
signal V_A_CTRL_LD_shadow_intermed_1 : STD_ULOGIC;
signal R_A_CTRL_INST19_intermed_2 : STD_LOGIC;
signal RIN_X_MEXC_intermed_1 : STD_ULOGIC;
signal RIN_D_MEXC_intermed_4 : STD_ULOGIC;
signal RIN_A_MULSTART_intermed_1 : STD_ULOGIC;
signal RIN_A_CTRL_TT_intermed_1 : std_logic_vector(5 downto 0);
signal RIN_M_CTRL_TT3DOWNTO0_intermed_2 : std_logic_vector(3 downto 0);
signal R_D_INST1_intermed_1 : std_logic_vector(31 downto 0);
signal RIN_A_CTRL_intermed_1 : PIPELINE_CTRL_TYPE;
signal R_E_CTRL_WICC_intermed_1 : STD_ULOGIC;
signal RIN_M_CTRL_TT3DOWNTO0_intermed_3 : std_logic_vector(3 downto 0);
signal V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 : std_logic_vector(31 downto 2);
signal V_A_CTRL_TT3DOWNTO0_shadow_intermed_1 : std_logic_vector(3 downto 0);
signal RIN_M_DCI_SIGNED_intermed_2 : STD_ULOGIC;
signal V_E_CTRL_TT3DOWNTO0_shadow_intermed_3 : std_logic_vector(3 downto 0);
signal IRIN_ADDR31DOWNTO4_intermed_1 : std_logic_vector(31 downto 4);
signal RIN_X_SET_intermed_1 : STD_LOGIC_VECTOR(0 downto 0);
signal V_M_CTRL_WREG_shadow_intermed_2 : STD_ULOGIC;
signal RIN_X_CTRL_PC31DOWNTO12_intermed_4 : std_logic_vector(31 downto 12);
signal V_D_PC_shadow_intermed_5 : std_logic_vector(31 downto 2);
signal RIN_X_CTRL_TT3DOWNTO0_intermed_2 : std_logic_vector(3 downto 0);
signal R_D_INST0_intermed_1 : std_logic_vector(31 downto 0);
signal R_E_CTRL_PC31DOWNTO4_intermed_4 : std_logic_vector(31 downto 4);
signal RIN_D_CNT_intermed_1 : std_logic_vector(1 downto 0);
signal R_E_CTRL_PC3DOWNTO2_intermed_4 : std_logic_vector(3 downto 2);
signal V_M_DCI_SIGNED_shadow_intermed_2 : STD_ULOGIC;
signal R_D_CNT_intermed_2 : std_logic_vector(1 downto 0);
signal R_E_CTRL_INST20_intermed_1 : STD_LOGIC;
signal RIN_M_DCI_SIGNED_intermed_1 : STD_ULOGIC;
signal RIN_D_PC3DOWNTO2_intermed_5 : std_logic_vector(3 downto 2);
signal RIN_A_CTRL_INST19_intermed_3 : STD_LOGIC;
signal V_E_CTRL_shadow_intermed_1 : PIPELINE_CTRL_TYPE;
signal RIN_A_CTRL_WICC_intermed_1 : STD_ULOGIC;
signal V_X_DATA1_shadow_intermed_1 : std_logic_vector(31 downto 0);
signal RIN_D_CWP_intermed_2 : std_logic_vector(2 downto 0);
signal R_E_CTRL_INST24_intermed_2 : STD_LOGIC;
signal V_A_CTRL_WREG_shadow_intermed_2 : STD_ULOGIC;
signal DCO_DATA031_intermed_2 : STD_LOGIC;
signal R_M_CTRL_TT_intermed_1 : std_logic_vector(5 downto 0);
signal RIN_E_CTRL_WREG_intermed_3 : STD_ULOGIC;
signal V_E_YMSB_shadow_intermed_1 : STD_ULOGIC;
signal IRIN_ADDR31DOWNTO2_intermed_3 : std_logic_vector(31 downto 2);
signal EX_JUMP_ADDRESS3DOWNTO2_shadow_intermed_1 : std_logic_vector(3 downto 2);
signal V_M_CTRL_INST_shadow_intermed_2 : std_logic_vector(31 downto 0);
signal DE_INST24_shadow_intermed_3 : STD_LOGIC;
signal V_D_PC31DOWNTO12_shadow_intermed_2 : std_logic_vector(31 downto 12);
signal V_A_CTRL_PC_shadow_intermed_1 : std_logic_vector(31 downto 2);
signal RIN_X_RESULT6DOWNTO0_intermed_1 : std_logic_vector(6 downto 0);
signal R_A_CTRL_PC31DOWNTO2_intermed_2 : std_logic_vector(31 downto 2);
signal V_E_CTRL_CNT_shadow_intermed_1 : std_logic_vector(1 downto 0);
signal VIR_ADDR3DOWNTO2_shadow_intermed_1 : std_logic_vector(3 downto 2);
signal RIN_A_CTRL_INST_intermed_2 : std_logic_vector(31 downto 0);
signal RIN_A_CTRL_intermed_3 : PIPELINE_CTRL_TYPE;
signal RIN_M_RESULT1DOWNTO0_intermed_1 : std_logic_vector(1 downto 0);
signal R_A_CTRL_PV_intermed_3 : STD_ULOGIC;
signal R_D_PC31DOWNTO2_intermed_1 : std_logic_vector(31 downto 2);
signal R_A_CTRL_PC31DOWNTO4_intermed_5 : std_logic_vector(31 downto 4);
signal RIN_A_DIVSTART_intermed_1 : STD_ULOGIC;
signal VIR_ADDR31DOWNTO12_shadow_intermed_2 : std_logic_vector(31 downto 12);
signal V_E_CTRL_INST20_shadow_intermed_2 : STD_LOGIC;
signal RIN_M_CTRL_TT_intermed_1 : std_logic_vector(5 downto 0);
signal RIN_E_CTRL_RD7DOWNTO0_intermed_3 : std_logic_vector(7 downto 0);
signal RIN_D_CWP_intermed_1 : std_logic_vector(2 downto 0);
signal RIN_X_CTRL_WREG_intermed_1 : STD_ULOGIC;
signal RIN_X_CTRL_PC31DOWNTO2_intermed_4 : std_logic_vector(31 downto 2);
signal V_M_CTRL_PC31DOWNTO2_shadow_intermed_5 : std_logic_vector(31 downto 2);
signal RIN_D_PC31DOWNTO2_intermed_7 : std_logic_vector(31 downto 2);
signal RIN_X_CTRL_PC31DOWNTO2_intermed_1 : std_logic_vector(31 downto 2);
signal DSUR_CRDY2_intermed_1 : STD_LOGIC;
signal R_E_CTRL_PC3DOWNTO2_intermed_2 : std_logic_vector(3 downto 2);
signal V_A_CTRL_RD7DOWNTO0_shadow_intermed_1 : std_logic_vector(7 downto 0);
signal R_D_PC31DOWNTO12_intermed_3 : std_logic_vector(31 downto 12);
signal RIN_X_DATA031_intermed_2 : STD_LOGIC;
signal RIN_D_PC31DOWNTO4_intermed_4 : std_logic_vector(31 downto 4);
signal RIN_A_CTRL_INST_intermed_4 : std_logic_vector(31 downto 0);
signal V_X_CTRL_PC31DOWNTO2_shadow_intermed_2 : std_logic_vector(31 downto 2);
signal V_M_CTRL_PC31DOWNTO4_shadow_intermed_2 : std_logic_vector(31 downto 4);
signal DE_INST19_shadow_intermed_1 : STD_LOGIC;
signal RIN_E_CTRL_PC31DOWNTO2_intermed_3 : std_logic_vector(31 downto 2);
signal V_A_CTRL_RD7DOWNTO0_shadow_intermed_2 : std_logic_vector(7 downto 0);
signal V_E_CTRL_INST_shadow_intermed_3 : std_logic_vector(31 downto 0);
signal RIN_X_CTRL_PC31DOWNTO2_intermed_2 : std_logic_vector(31 downto 2);
signal RIN_X_CTRL_intermed_1 : PIPELINE_CTRL_TYPE;
signal R_D_PC31DOWNTO12_intermed_1 : std_logic_vector(31 downto 12);
signal RIN_A_CTRL_ANNUL_intermed_2 : STD_ULOGIC;
signal V_A_CTRL_CNT_shadow_intermed_3 : std_logic_vector(1 downto 0);
signal R_A_CTRL_PC31DOWNTO12_intermed_6 : std_logic_vector(31 downto 12);
signal V_M_CTRL_PC31DOWNTO12_shadow_intermed_4 : std_logic_vector(31 downto 12);
signal VIR_ADDR31DOWNTO2_shadow_intermed_3 : std_logic_vector(31 downto 2);
signal V_A_MULSTART_shadow_intermed_1 : STD_ULOGIC;
signal RIN_X_DATA1_intermed_2 : std_logic_vector(31 downto 0);
signal RIN_E_CTRL_PC_intermed_2 : std_logic_vector(31 downto 2);
signal V_E_CTRL_PC31DOWNTO12_shadow_intermed_5 : std_logic_vector(31 downto 12);
signal V_M_DCI_SIZE_shadow_intermed_1 : std_logic_vector(1 downto 0);
signal V_A_CTRL_PC31DOWNTO4_shadow_intermed_3 : std_logic_vector(31 downto 4);
signal R_X_RESULT6DOWNTO03DOWNTO0_intermed_3 : std_logic_vector(3 downto 0);
signal R_D_PC31DOWNTO4_intermed_6 : std_logic_vector(31 downto 4);
signal EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_2 : STD_LOGIC_VECTOR(32 downto 3);
signal V_A_CTRL_PV_shadow_intermed_4 : STD_ULOGIC;
signal V_A_CTRL_TT_shadow_intermed_4 : std_logic_vector(5 downto 0);
signal V_X_CTRL_PC3DOWNTO2_shadow_intermed_3 : std_logic_vector(3 downto 2);
signal RIN_X_DATA0_intermed_2 : std_logic_vector(31 downto 0);
signal R_A_CTRL_TT3DOWNTO0_intermed_4 : std_logic_vector(3 downto 0);
signal RIN_D_PC31DOWNTO4_intermed_3 : std_logic_vector(31 downto 4);
signal V_A_CTRL_WREG_shadow_intermed_4 : STD_ULOGIC;
signal RIN_A_CTRL_PC3DOWNTO2_intermed_1 : std_logic_vector(3 downto 2);
signal RIN_D_PC31DOWNTO2_intermed_2 : std_logic_vector(31 downto 2);
signal R_M_CTRL_PC_intermed_2 : std_logic_vector(31 downto 2);
signal R_F_PC31DOWNTO2_intermed_2 : std_logic_vector(31 downto 2);
signal RIN_M_CTRL_WREG_intermed_1 : STD_ULOGIC;
signal RIN_W_WREG_intermed_1 : STD_ULOGIC;
signal RIN_D_PC31DOWNTO4_intermed_6 : std_logic_vector(31 downto 4);
signal R_D_ANNUL_intermed_1 : STD_ULOGIC;
signal R_A_CTRL_INST_intermed_3 : std_logic_vector(31 downto 0);
signal RIN_M_CTRL_PC31DOWNTO2_intermed_2 : std_logic_vector(31 downto 2);
signal RIN_E_CTRL_WREG_intermed_2 : STD_ULOGIC;
signal V_E_SARI_shadow_intermed_1 : STD_ULOGIC;
signal R_E_CTRL_RD6DOWNTO0_intermed_2 : std_logic_vector(6 downto 0);
signal V_A_CTRL_PC31DOWNTO2_shadow_intermed_6 : std_logic_vector(31 downto 2);
signal R_A_CTRL_CNT_intermed_3 : std_logic_vector(1 downto 0);
signal RIN_M_CTRL_PV_intermed_2 : STD_ULOGIC;
signal R_A_CTRL_LD_intermed_1 : STD_ULOGIC;
signal V_E_CTRL_WICC_shadow_intermed_2 : STD_ULOGIC;
signal RIN_D_PC31DOWNTO2_intermed_5 : std_logic_vector(31 downto 2);
signal V_D_PC3DOWNTO2_shadow_intermed_3 : std_logic_vector(3 downto 2);
signal RIN_A_CTRL_PC3DOWNTO2_intermed_6 : std_logic_vector(3 downto 2);
signal RIN_X_DATA04DOWNTO0_intermed_1 : std_logic_vector(4 downto 0);
signal DSUIN_CRDY2_intermed_1 : STD_LOGIC;
signal RIN_D_PC31DOWNTO12_intermed_4 : std_logic_vector(31 downto 12);
signal R_E_CTRL_RD6DOWNTO0_intermed_1 : std_logic_vector(6 downto 0);
signal RIN_A_CTRL_INST20_intermed_1 : STD_LOGIC;
signal R_M_RESULT1DOWNTO0_intermed_2 : std_logic_vector(1 downto 0);
signal RIN_M_DCI_SIZE_intermed_2 : std_logic_vector(1 downto 0);
signal DE_INST19_shadow_intermed_3 : STD_LOGIC;
signal IRIN_ADDR31DOWNTO12_intermed_2 : std_logic_vector(31 downto 12);
signal V_A_CTRL_ANNUL_shadow_intermed_4 : STD_ULOGIC;
signal R_E_CTRL_CNT_intermed_1 : std_logic_vector(1 downto 0);
signal V_E_CTRL_INST24_shadow_intermed_2 : STD_LOGIC;
signal RIN_A_CTRL_PC31DOWNTO4_intermed_2 : std_logic_vector(31 downto 4);
signal IRIN_PWD_intermed_1 : STD_ULOGIC;
signal V_D_MEXC_shadow_intermed_5 : STD_ULOGIC;
signal RIN_A_CTRL_PV_intermed_1 : STD_ULOGIC;
signal V_A_CTRL_WICC_shadow_intermed_1 : STD_ULOGIC;
signal R_A_CTRL_PC_intermed_1 : std_logic_vector(31 downto 2);
signal V_F_PC31DOWNTO4_shadow_intermed_1 : std_logic_vector(31 downto 4);
signal R_A_CTRL_RD7DOWNTO0_intermed_3 : std_logic_vector(7 downto 0);
signal RIN_A_CTRL_PC_intermed_1 : std_logic_vector(31 downto 2);
signal R_E_CTRL_INST_intermed_1 : std_logic_vector(31 downto 0);
signal R_E_CTRL_PC31DOWNTO4_intermed_1 : std_logic_vector(31 downto 4);
signal V_A_CTRL_TRAP_shadow_intermed_4 : STD_ULOGIC;
signal V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 : std_logic_vector(31 downto 2);
signal V_F_PC31DOWNTO12_shadow_intermed_1 : std_logic_vector(31 downto 12);
signal R_A_CTRL_PC3DOWNTO2_intermed_5 : std_logic_vector(3 downto 2);
signal R_A_CTRL_CNT_intermed_1 : std_logic_vector(1 downto 0);
signal RIN_D_PC31DOWNTO2_intermed_6 : std_logic_vector(31 downto 2);
signal R_E_CTRL_PC3DOWNTO2_intermed_1 : std_logic_vector(3 downto 2);
signal RIN_X_DATA0_intermed_1 : std_logic_vector(31 downto 0);
signal RIN_E_CTRL_PC_intermed_3 : std_logic_vector(31 downto 2);
signal R_X_CTRL_PC31DOWNTO12_intermed_1 : std_logic_vector(31 downto 12);
signal RIN_X_DATA03_intermed_1 : STD_LOGIC;
signal R_X_DATA04DOWNTO0_intermed_2 : std_logic_vector(4 downto 0);
signal R_E_CTRL_ANNUL_intermed_1 : STD_ULOGIC;
signal V_A_CTRL_RD7DOWNTO0_shadow_intermed_3 : std_logic_vector(7 downto 0);
signal V_M_CTRL_TT3DOWNTO0_shadow_intermed_3 : std_logic_vector(3 downto 0);
signal RIN_X_MAC_intermed_1 : STD_ULOGIC;
signal V_E_SHCNT_shadow_intermed_1 : std_logic_vector(4 downto 0);
signal V_M_CTRL_TT3DOWNTO0_shadow_intermed_2 : std_logic_vector(3 downto 0);
signal V_D_PC31DOWNTO12_shadow_intermed_4 : std_logic_vector(31 downto 12);
signal RIN_D_PC31DOWNTO12_intermed_2 : std_logic_vector(31 downto 12);
signal V_E_CTRL_PC3DOWNTO2_shadow_intermed_5 : std_logic_vector(3 downto 2);
signal RIN_E_CTRL_RETT_intermed_2 : STD_ULOGIC;
signal R_M_CTRL_PC31DOWNTO2_intermed_2 : std_logic_vector(31 downto 2);
signal V_E_OP23_shadow_intermed_1 : STD_LOGIC;
signal V_D_PC_shadow_intermed_2 : std_logic_vector(31 downto 2);
signal R_D_PC3DOWNTO2_intermed_6 : std_logic_vector(3 downto 2);
signal R_M_CTRL_PV_intermed_1 : STD_ULOGIC;
signal RIN_W_RESULT_intermed_1 : std_logic_vector(31 downto 0);
signal V_E_CTRL_ANNUL_shadow_intermed_2 : STD_ULOGIC;
signal V_E_CTRL_PV_shadow_intermed_1 : STD_ULOGIC;
signal RIN_X_LADDR_intermed_1 : std_logic_vector(1 downto 0);
signal RIN_A_CTRL_PC_intermed_5 : std_logic_vector(31 downto 2);
signal XC_VECTT3DOWNTO0_shadow_intermed_1 : STD_LOGIC_VECTOR(3 downto 0);
signal R_E_CTRL_WREG_intermed_1 : STD_ULOGIC;
signal RIN_X_DATA03_intermed_2 : STD_LOGIC;
signal RIN_A_CTRL_TT_intermed_3 : std_logic_vector(5 downto 0);
signal V_D_STEP_shadow_intermed_1 : STD_ULOGIC;
signal R_M_CTRL_PC31DOWNTO12_intermed_1 : std_logic_vector(31 downto 12);
signal DE_INST19_shadow_intermed_2 : STD_LOGIC;
signal RIN_M_CTRL_PC31DOWNTO2_intermed_3 : std_logic_vector(31 downto 2);
signal V_X_CTRL_TRAP_shadow_intermed_1 : STD_ULOGIC;
signal RIN_D_MEXC_intermed_5 : STD_ULOGIC;
signal RIN_X_CTRL_TRAP_intermed_1 : STD_ULOGIC;
signal V_D_PC3DOWNTO2_shadow_intermed_4 : std_logic_vector(3 downto 2);
signal V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1 : std_logic_vector(3 downto 0);
signal RIN_A_CTRL_PC3DOWNTO2_intermed_5 : std_logic_vector(3 downto 2);
signal RIN_M_CTRL_PC31DOWNTO4_intermed_3 : std_logic_vector(31 downto 4);
signal RIN_M_CTRL_PC31DOWNTO2_intermed_4 : std_logic_vector(31 downto 2);
signal RIN_F_BRANCH_intermed_1 : STD_ULOGIC;
signal R_D_PC3DOWNTO2_intermed_5 : std_logic_vector(3 downto 2);
signal RIN_A_CTRL_WREG_intermed_1 : STD_ULOGIC;
signal RIN_D_INST0_intermed_2 : std_logic_vector(31 downto 0);
signal R_M_CTRL_CNT_intermed_1 : std_logic_vector(1 downto 0);
signal RIN_E_CTRL_RD7DOWNTO0_intermed_1 : std_logic_vector(7 downto 0);
signal RIN_A_CTRL_PC_intermed_2 : std_logic_vector(31 downto 2);
signal RIN_X_CTRL_PC_intermed_1 : std_logic_vector(31 downto 2);
signal R_A_SU_intermed_1 : STD_ULOGIC;
signal RIN_A_CTRL_TT_intermed_4 : std_logic_vector(5 downto 0);
signal V_X_DATA00_shadow_intermed_2 : STD_LOGIC;
signal RIN_A_CTRL_PC31DOWNTO4_intermed_4 : std_logic_vector(31 downto 4);
signal RIN_A_JMPL_intermed_1 : STD_ULOGIC;
signal V_E_CTRL_WREG_shadow_intermed_3 : STD_ULOGIC;
signal V_A_CTRL_WREG_shadow_intermed_1 : STD_ULOGIC;
signal RIN_M_CTRL_ANNUL_intermed_1 : STD_ULOGIC;
signal RIN_X_CTRL_PC31DOWNTO12_intermed_1 : std_logic_vector(31 downto 12);
signal VIR_ADDR31DOWNTO2_shadow_intermed_1 : std_logic_vector(31 downto 2);
signal V_A_CTRL_PC3DOWNTO2_shadow_intermed_1 : std_logic_vector(3 downto 2);
signal RIN_E_CTRL_TT3DOWNTO0_intermed_3 : std_logic_vector(3 downto 0);
signal RIN_M_CTRL_RD7DOWNTO0_intermed_2 : std_logic_vector(7 downto 0);
signal V_E_CTRL_TRAP_shadow_intermed_3 : STD_ULOGIC;
signal V_A_CTRL_CNT_shadow_intermed_2 : std_logic_vector(1 downto 0);
signal V_E_CTRL_ANNUL_shadow_intermed_1 : STD_ULOGIC;
signal V_W_S_TT3DOWNTO0_shadow_intermed_1 : STD_LOGIC_VECTOR(3 downto 0);
signal RIN_M_CTRL_CNT_intermed_1 : std_logic_vector(1 downto 0);
signal DSUR_CRDY2_intermed_2 : STD_LOGIC;
signal V_E_CTRL_RD6DOWNTO0_shadow_intermed_1 : std_logic_vector(6 downto 0);
signal V_A_CTRL_CNT_shadow_intermed_1 : std_logic_vector(1 downto 0);
signal R_E_CTRL_PC_intermed_1 : std_logic_vector(31 downto 2);
signal RIN_M_SU_intermed_1 : STD_ULOGIC;
signal RIN_A_CTRL_RD6DOWNTO0_intermed_1 : std_logic_vector(6 downto 0);
signal R_M_CTRL_TT3DOWNTO0_intermed_3 : std_logic_vector(3 downto 0);
signal RIN_M_CTRL_TT3DOWNTO0_intermed_4 : std_logic_vector(3 downto 0);
signal V_A_CTRL_INST19_shadow_intermed_1 : STD_LOGIC;
signal R_D_PC31DOWNTO2_intermed_5 : std_logic_vector(31 downto 2);
signal RIN_E_CTRL_CNT_intermed_3 : std_logic_vector(1 downto 0);
signal R_E_CTRL_PC31DOWNTO12_intermed_3 : std_logic_vector(31 downto 12);
signal RIN_E_CTRL_TRAP_intermed_1 : STD_ULOGIC;
signal RIN_X_DATA00_intermed_3 : STD_LOGIC;
signal R_E_CTRL_PC_intermed_2 : std_logic_vector(31 downto 2);
signal RIN_E_OP131_intermed_1 : STD_LOGIC;
signal R_D_CNT_intermed_1 : std_logic_vector(1 downto 0);
signal R_D_PC_intermed_3 : std_logic_vector(31 downto 2);
signal RIN_A_CTRL_PC31DOWNTO12_intermed_2 : std_logic_vector(31 downto 12);
signal R_M_CTRL_WREG_intermed_1 : STD_ULOGIC;
signal R_D_PC31DOWNTO2_intermed_4 : std_logic_vector(31 downto 2);
signal DE_INST_shadow_intermed_3 : std_logic_vector(31 downto 0);
signal RIN_D_PC_intermed_3 : std_logic_vector(31 downto 2);
signal V_A_CTRL_INST20_shadow_intermed_3 : STD_LOGIC;
signal R_A_CTRL_TT3DOWNTO0_intermed_5 : std_logic_vector(3 downto 0);
signal RIN_A_CTRL_CNT_intermed_2 : std_logic_vector(1 downto 0);
signal RIN_A_CTRL_intermed_2 : PIPELINE_CTRL_TYPE;
signal RIN_X_CTRL_PC_intermed_2 : std_logic_vector(31 downto 2);
signal R_A_CTRL_WREG_intermed_1 : STD_ULOGIC;
signal V_X_CTRL_PC31DOWNTO2_shadow_intermed_4 : std_logic_vector(31 downto 2);
signal R_X_CTRL_PC31DOWNTO2_intermed_3 : std_logic_vector(31 downto 2);
signal RIN_D_PC_intermed_6 : std_logic_vector(31 downto 2);
signal RIN_E_CTRL_PC31DOWNTO4_intermed_3 : std_logic_vector(31 downto 4);
signal R_X_CTRL_PC31DOWNTO2_intermed_2 : std_logic_vector(31 downto 2);
signal V_A_ET_shadow_intermed_1 : STD_ULOGIC;
signal V_E_CTRL_PC31DOWNTO4_shadow_intermed_1 : std_logic_vector(31 downto 4);
signal RIN_A_CTRL_INST20_intermed_3 : STD_LOGIC;
signal RIN_W_EXCEPT_intermed_1 : STD_ULOGIC;
signal V_X_DATA031_shadow_intermed_2 : STD_LOGIC;
signal R_A_CTRL_ANNUL_intermed_1 : STD_ULOGIC;
signal R_F_PC31DOWNTO12_intermed_1 : std_logic_vector(31 downto 12);
signal RIN_E_CTRL_RD6DOWNTO0_intermed_2 : std_logic_vector(6 downto 0);
signal VIR_ADDR31DOWNTO2_shadow_intermed_2 : std_logic_vector(31 downto 2);
signal RIN_X_DATA00_intermed_1 : STD_LOGIC;
signal RIN_E_CTRL_ANNUL_intermed_1 : STD_ULOGIC;
signal RIN_E_CTRL_PC31DOWNTO4_intermed_5 : std_logic_vector(31 downto 4);
signal V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_3 : std_logic_vector(3 downto 0);
signal V_M_CTRL_WICC_shadow_intermed_1 : STD_ULOGIC;
signal V_A_CTRL_PC31DOWNTO2_shadow_intermed_7 : std_logic_vector(31 downto 2);
signal RIN_A_CTRL_RETT_intermed_1 : STD_ULOGIC;
signal RIN_E_CTRL_PC31DOWNTO2_intermed_1 : std_logic_vector(31 downto 2);
signal V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 : std_logic_vector(31 downto 2);
signal RIN_D_PC31DOWNTO12_intermed_5 : std_logic_vector(31 downto 12);
signal VIR_ADDR3DOWNTO2_shadow_intermed_2 : std_logic_vector(3 downto 2);
signal R_A_CTRL_PV_intermed_2 : STD_ULOGIC;
signal V_A_CTRL_PC3DOWNTO2_shadow_intermed_2 : std_logic_vector(3 downto 2);
signal R_E_CTRL_PC3DOWNTO2_intermed_3 : std_logic_vector(3 downto 2);
signal V_A_CTRL_ANNUL_shadow_intermed_3 : STD_ULOGIC;
signal RIN_A_CTRL_PC3DOWNTO2_intermed_4 : std_logic_vector(3 downto 2);
signal V_A_CTRL_TT3DOWNTO0_shadow_intermed_3 : std_logic_vector(3 downto 0);
signal R_A_CTRL_PC3DOWNTO2_intermed_2 : std_logic_vector(3 downto 2);
signal V_D_CNT_shadow_intermed_2 : std_logic_vector(1 downto 0);
signal V_M_CTRL_ANNUL_shadow_intermed_1 : STD_ULOGIC;
signal V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 : std_logic_vector(31 downto 2);
signal RIN_M_CTRL_PC31DOWNTO4_intermed_2 : std_logic_vector(31 downto 4);
signal R_M_CTRL_TT3DOWNTO0_intermed_1 : std_logic_vector(3 downto 0);
signal V_E_CTRL_LD_shadow_intermed_2 : STD_ULOGIC;
signal RIN_X_CTRL_ANNUL_intermed_1 : STD_ULOGIC;
signal RIN_D_PC3DOWNTO2_intermed_3 : std_logic_vector(3 downto 2);
signal V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 : std_logic_vector(31 downto 2);
signal RIN_E_CTRL_TT_intermed_2 : std_logic_vector(5 downto 0);
signal RIN_E_CTRL_CNT_intermed_2 : std_logic_vector(1 downto 0);
signal RIN_A_CTRL_PC_intermed_4 : std_logic_vector(31 downto 2);
signal RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_4 : std_logic_vector(3 downto 0);
signal R_D_PC31DOWNTO12_intermed_2 : std_logic_vector(31 downto 12);
signal XC_TRAP_ADDRESS31DOWNTO4_shadow_intermed_1 : std_logic_vector(31 downto 4);
signal RIN_A_CTRL_INST24_intermed_3 : STD_LOGIC;
signal V_W_S_TT3DOWNTO0_shadow_intermed_2 : STD_LOGIC_VECTOR(3 downto 0);
signal RIN_E_CTRL_RD7DOWNTO0_intermed_2 : std_logic_vector(7 downto 0);
signal RIN_A_CTRL_INST24_intermed_1 : STD_LOGIC;
signal RIN_D_PC31DOWNTO4_intermed_2 : std_logic_vector(31 downto 4);
signal V_A_CTRL_shadow_intermed_2 : PIPELINE_CTRL_TYPE;
signal DE_INST_shadow_intermed_4 : std_logic_vector(31 downto 0);
signal RIN_E_CTRL_PV_intermed_3 : STD_ULOGIC;
signal V_A_CTRL_TT_shadow_intermed_2 : std_logic_vector(5 downto 0);
signal RIN_M_CTRL_PC_intermed_3 : std_logic_vector(31 downto 2);
signal V_A_CTRL_WREG_shadow_intermed_3 : STD_ULOGIC;
signal R_M_CTRL_RD6DOWNTO0_intermed_1 : std_logic_vector(6 downto 0);
signal XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_1 : std_logic_vector(31 downto 2);
signal RIN_A_CTRL_PV_intermed_2 : STD_ULOGIC;
signal RIN_E_CTRL_PC3DOWNTO2_intermed_2 : std_logic_vector(3 downto 2);
signal RIN_X_CTRL_RD7DOWNTO0_intermed_1 : std_logic_vector(7 downto 0);
signal V_A_CTRL_TRAP_shadow_intermed_1 : STD_ULOGIC;
signal V_E_CTRL_TRAP_shadow_intermed_1 : STD_ULOGIC;
signal RIN_E_MAC_intermed_1 : STD_ULOGIC;
signal R_X_DATA00_intermed_2 : STD_LOGIC;
signal RIN_E_MAC_intermed_2 : STD_ULOGIC;
signal RIN_A_CTRL_RD7DOWNTO0_intermed_4 : std_logic_vector(7 downto 0);
signal RIN_A_CTRL_PC31DOWNTO2_intermed_7 : std_logic_vector(31 downto 2);
signal R_M_CTRL_PC31DOWNTO12_intermed_3 : std_logic_vector(31 downto 12);
signal V_D_PC_shadow_intermed_3 : std_logic_vector(31 downto 2);
signal RIN_D_PC31DOWNTO4_intermed_5 : std_logic_vector(31 downto 4);
signal V_M_RESULT1DOWNTO0_shadow_intermed_2 : std_logic_vector(1 downto 0);
signal R_E_CTRL_PC31DOWNTO4_intermed_2 : std_logic_vector(31 downto 4);
signal V_E_CTRL_PC31DOWNTO12_shadow_intermed_3 : std_logic_vector(31 downto 12);
signal V_X_INTACK_shadow_intermed_1 : STD_ULOGIC;
signal RIN_A_CTRL_ANNUL_intermed_5 : STD_ULOGIC;
signal V_M_CTRL_PC31DOWNTO4_shadow_intermed_3 : std_logic_vector(31 downto 4);
signal V_A_CTRL_TT3DOWNTO0_shadow_intermed_4 : std_logic_vector(3 downto 0);
signal RIN_X_RESULT_intermed_1 : std_logic_vector(31 downto 0);
signal RIN_E_CTRL_TT3DOWNTO0_intermed_5 : std_logic_vector(3 downto 0);
signal RIN_A_CTRL_PC31DOWNTO2_intermed_1 : std_logic_vector(31 downto 2);
signal EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_1 : std_logic_vector(31 downto 2);
signal V_D_PC3DOWNTO2_shadow_intermed_5 : std_logic_vector(3 downto 2);
signal DE_INST20_shadow_intermed_1 : STD_LOGIC;
signal V_E_CTRL_RD7DOWNTO0_shadow_intermed_2 : std_logic_vector(7 downto 0);
signal V_X_CTRL_PC31DOWNTO12_shadow_intermed_4 : std_logic_vector(31 downto 12);
signal V_E_CTRL_TRAP_shadow_intermed_2 : STD_ULOGIC;
signal V_A_CTRL_PC31DOWNTO4_shadow_intermed_5 : std_logic_vector(31 downto 4);
signal V_A_CTRL_RD6DOWNTO0_shadow_intermed_2 : std_logic_vector(6 downto 0);
signal RIN_A_CTRL_PC31DOWNTO12_intermed_1 : std_logic_vector(31 downto 12);
signal IR_ADDR31DOWNTO12_intermed_2 : std_logic_vector(31 downto 12);
signal RIN_E_ALUCIN_intermed_1 : STD_ULOGIC;
signal R_X_CTRL_PC31DOWNTO12_intermed_2 : std_logic_vector(31 downto 12);
signal R_A_CTRL_PC3DOWNTO2_intermed_1 : std_logic_vector(3 downto 2);
signal DE_INST_shadow_intermed_1 : std_logic_vector(31 downto 0);
signal RIN_M_CTRL_INST_intermed_2 : std_logic_vector(31 downto 0);
signal R_A_CTRL_TRAP_intermed_2 : STD_ULOGIC;
signal RIN_A_CTRL_PC31DOWNTO12_intermed_4 : std_logic_vector(31 downto 12);
signal R_A_CTRL_WREG_intermed_2 : STD_ULOGIC;
signal R_M_CTRL_PC31DOWNTO4_intermed_1 : std_logic_vector(31 downto 4);
signal V_E_OP13_shadow_intermed_1 : STD_LOGIC;
signal V_A_CTRL_INST24_shadow_intermed_1 : STD_LOGIC;
signal V_X_CTRL_PC31DOWNTO12_shadow_intermed_3 : std_logic_vector(31 downto 12);
signal IRIN_ADDR31DOWNTO12_intermed_3 : std_logic_vector(31 downto 12);
signal V_X_CTRL_PC_shadow_intermed_1 : std_logic_vector(31 downto 2);
signal R_M_CTRL_PC3DOWNTO2_intermed_3 : std_logic_vector(3 downto 2);
signal V_E_CTRL_PC3DOWNTO2_shadow_intermed_2 : std_logic_vector(3 downto 2);
signal RIN_X_CTRL_TT_intermed_1 : std_logic_vector(5 downto 0);
signal V_M_CTRL_PC31DOWNTO2_shadow_intermed_3 : std_logic_vector(31 downto 2);
signal RIN_A_CTRL_TT3DOWNTO0_intermed_6 : std_logic_vector(3 downto 0);
signal RIN_D_PC3DOWNTO2_intermed_7 : std_logic_vector(3 downto 2);
signal V_A_CTRL_INST_shadow_intermed_2 : std_logic_vector(31 downto 0);
signal V_X_CTRL_PC31DOWNTO4_shadow_intermed_1 : std_logic_vector(31 downto 4);
signal V_M_RESULT1DOWNTO0_shadow_intermed_1 : std_logic_vector(1 downto 0);
signal R_A_CTRL_INST24_intermed_2 : STD_LOGIC;
signal R_F_PC31DOWNTO2_intermed_1 : std_logic_vector(31 downto 2);
signal V_A_CTRL_TRAP_shadow_intermed_3 : STD_ULOGIC;
signal R_D_CNT_intermed_4 : std_logic_vector(1 downto 0);
signal RIN_A_CTRL_WREG_intermed_4 : STD_ULOGIC;
signal V_M_CTRL_PC31DOWNTO4_shadow_intermed_1 : std_logic_vector(31 downto 4);
signal RIN_A_CTRL_PC3DOWNTO2_intermed_3 : std_logic_vector(3 downto 2);
signal V_E_CTRL_INST20_shadow_intermed_1 : STD_LOGIC;
signal R_D_MEXC_intermed_2 : STD_ULOGIC;
signal R_D_PC_intermed_4 : std_logic_vector(31 downto 2);
signal RIN_D_PC_intermed_1 : std_logic_vector(31 downto 2);
signal IRIN_ADDR3DOWNTO2_intermed_1 : std_logic_vector(3 downto 2);
signal V_E_CTRL_RD7DOWNTO0_shadow_intermed_1 : std_logic_vector(7 downto 0);
signal RIN_E_OP1_intermed_1 : std_logic_vector(31 downto 0);
signal V_D_PC31DOWNTO4_shadow_intermed_3 : std_logic_vector(31 downto 4);
signal V_A_CTRL_PV_shadow_intermed_3 : STD_ULOGIC;
signal V_D_PC31DOWNTO2_shadow_intermed_6 : std_logic_vector(31 downto 2);
signal V_X_CTRL_TT3DOWNTO0_shadow_intermed_2 : std_logic_vector(3 downto 0);
signal DE_INST20_shadow_intermed_2 : STD_LOGIC;
signal V_E_CTRL_RD7DOWNTO0_shadow_intermed_3 : std_logic_vector(7 downto 0);
signal V_E_CTRL_CNT_shadow_intermed_3 : std_logic_vector(1 downto 0);
signal RIN_E_CTRL_RETT_intermed_1 : STD_ULOGIC;
signal V_D_PC31DOWNTO12_shadow_intermed_3 : std_logic_vector(31 downto 12);
signal V_D_PC31DOWNTO12_shadow_intermed_7 : std_logic_vector(31 downto 12);
signal V_M_CTRL_CNT_shadow_intermed_2 : std_logic_vector(1 downto 0);
signal R_D_PC31DOWNTO4_intermed_3 : std_logic_vector(31 downto 4);
signal RIN_A_CTRL_PC3DOWNTO2_intermed_2 : std_logic_vector(3 downto 2);
signal RIN_X_INTACK_intermed_1 : STD_ULOGIC;
signal RIN_E_OP231_intermed_1 : STD_LOGIC;
signal RIN_X_DATA031_intermed_3 : STD_LOGIC;
signal RIN_D_PC31DOWNTO2_intermed_4 : std_logic_vector(31 downto 2);
signal V_D_PC31DOWNTO4_shadow_intermed_2 : std_logic_vector(31 downto 4);
signal V_A_CTRL_ANNUL_shadow_intermed_1 : STD_ULOGIC;
signal R_M_CTRL_TT3DOWNTO0_intermed_2 : std_logic_vector(3 downto 0);
signal V_F_PC_shadow_intermed_1 : std_logic_vector(31 downto 2);
signal RIN_E_ET_intermed_1 : STD_ULOGIC;
signal V_D_MEXC_shadow_intermed_3 : STD_ULOGIC;
signal XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_2 : std_logic_vector(31 downto 2);
signal V_F_PC31DOWNTO2_shadow_intermed_2 : std_logic_vector(31 downto 2);
signal RIN_E_CTRL_PV_intermed_2 : STD_ULOGIC;
signal R_A_CTRL_RD7DOWNTO0_intermed_1 : std_logic_vector(7 downto 0);
signal ICO_MEXC_intermed_2 : STD_ULOGIC;
signal V_X_DCI_SIGNED_shadow_intermed_1 : STD_ULOGIC;
signal RIN_A_STEP_intermed_1 : STD_ULOGIC;
signal V_E_ALUCIN_shadow_intermed_1 : STD_ULOGIC;
signal V_A_CTRL_PC31DOWNTO4_shadow_intermed_6 : std_logic_vector(31 downto 4);
signal V_D_CNT_shadow_intermed_3 : std_logic_vector(1 downto 0);
signal V_D_PC31DOWNTO4_shadow_intermed_1 : std_logic_vector(31 downto 4);
signal RIN_X_CTRL_CNT_intermed_1 : std_logic_vector(1 downto 0);
signal V_D_ANNUL_shadow_intermed_1 : STD_ULOGIC;
signal V_E_CTRL_PC31DOWNTO2_shadow_intermed_5 : std_logic_vector(31 downto 2);
signal V_E_CTRL_PV_shadow_intermed_3 : STD_ULOGIC;
signal VP_ERROR_shadow_intermed_1 : STD_ULOGIC;
signal RIN_X_RESULT6DOWNTO0_intermed_2 : std_logic_vector(6 downto 0);
signal R_D_PC31DOWNTO4_intermed_1 : std_logic_vector(31 downto 4);
signal RIN_F_PC31DOWNTO2_intermed_1 : std_logic_vector(31 downto 2);
signal RIN_E_CTRL_PC_intermed_1 : std_logic_vector(31 downto 2);
signal R_A_CTRL_PC31DOWNTO12_intermed_1 : std_logic_vector(31 downto 12);
signal RIN_A_CTRL_PC31DOWNTO12_intermed_6 : std_logic_vector(31 downto 12);
signal V_A_CTRL_INST24_shadow_intermed_3 : STD_LOGIC;
signal V_E_CTRL_PC_shadow_intermed_1 : std_logic_vector(31 downto 2);
signal V_X_CTRL_RD7DOWNTO0_shadow_intermed_1 : std_logic_vector(7 downto 0);
signal RIN_M_MUL_intermed_1 : STD_ULOGIC;
signal RIN_A_CTRL_INST20_intermed_2 : STD_LOGIC;
signal RIN_A_CTRL_RD7DOWNTO0_intermed_1 : std_logic_vector(7 downto 0);
signal V_A_CTRL_TT3DOWNTO0_shadow_intermed_2 : std_logic_vector(3 downto 0);
signal R_A_CTRL_INST_intermed_2 : std_logic_vector(31 downto 0);
signal RIN_E_CTRL_PC31DOWNTO2_intermed_6 : std_logic_vector(31 downto 2);
signal V_M_CTRL_TT_shadow_intermed_2 : std_logic_vector(5 downto 0);
signal V_D_INST0_shadow_intermed_2 : std_logic_vector(31 downto 0);
signal DCO_DATA03_intermed_1 : STD_LOGIC;
signal RIN_M_CTRL_intermed_1 : PIPELINE_CTRL_TYPE;
signal RIN_A_CTRL_RD7DOWNTO0_intermed_3 : std_logic_vector(7 downto 0);
signal V_D_PC31DOWNTO2_shadow_intermed_1 : std_logic_vector(31 downto 2);
signal RIN_E_CTRL_PC31DOWNTO4_intermed_2 : std_logic_vector(31 downto 4);
signal V_D_PC31DOWNTO12_shadow_intermed_8 : std_logic_vector(31 downto 12);
signal RIN_E_CTRL_LD_intermed_1 : STD_ULOGIC;
signal R_X_CTRL_PC_intermed_1 : std_logic_vector(31 downto 2);
signal RIN_A_CTRL_WY_intermed_1 : STD_ULOGIC;
signal RIN_D_PC3DOWNTO2_intermed_1 : std_logic_vector(3 downto 2);
signal R_E_CTRL_INST24_intermed_1 : STD_LOGIC;
signal V_M_DCI_shadow_intermed_1 : DC_IN_TYPE;
signal V_M_CTRL_shadow_intermed_1 : PIPELINE_CTRL_TYPE;
signal RIN_M_DCI_SIZE_intermed_1 : std_logic_vector(1 downto 0);
signal R_E_CTRL_PV_intermed_2 : STD_ULOGIC;
signal EX_ADD_RES32DOWNTO3_shadow_intermed_1 : STD_LOGIC_VECTOR(32 downto 3);
signal RIN_D_MEXC_intermed_1 : STD_ULOGIC;
signal R_A_CTRL_PC31DOWNTO2_intermed_3 : std_logic_vector(31 downto 2);
signal DSUIN_TBUFCNT_intermed_1 : STD_LOGIC_VECTOR(6 downto 0);
signal R_E_CTRL_PC31DOWNTO12_intermed_5 : std_logic_vector(31 downto 12);
signal R_A_CTRL_PC3DOWNTO2_intermed_4 : std_logic_vector(3 downto 2);
signal V_A_CTRL_INST20_shadow_intermed_1 : STD_LOGIC;
signal RIN_E_CTRL_PC31DOWNTO12_intermed_3 : std_logic_vector(31 downto 12);
signal V_A_CTRL_RD6DOWNTO0_shadow_intermed_4 : std_logic_vector(6 downto 0);
signal R_E_CTRL_PC31DOWNTO2_intermed_4 : std_logic_vector(31 downto 2);
signal R_A_CTRL_TT3DOWNTO0_intermed_2 : std_logic_vector(3 downto 0);
signal RIN_A_CTRL_CNT_intermed_4 : std_logic_vector(1 downto 0);
signal V_D_INST1_shadow_intermed_2 : std_logic_vector(31 downto 0);
signal RIN_E_CTRL_INST_intermed_1 : std_logic_vector(31 downto 0);
signal RIN_X_DEBUG_intermed_1 : STD_ULOGIC;
signal RIN_M_Y_intermed_1 : std_logic_vector(31 downto 0);
signal RIN_E_SHCNT_intermed_1 : std_logic_vector(4 downto 0);
signal RIN_E_CTRL_TRAP_intermed_2 : STD_ULOGIC;
signal RIN_F_PC31DOWNTO12_intermed_2 : std_logic_vector(31 downto 12);
signal R_E_CTRL_INST20_intermed_2 : STD_LOGIC;
signal RIN_A_CTRL_ANNUL_intermed_3 : STD_ULOGIC;
signal RIN_D_ANNUL_intermed_2 : STD_ULOGIC;
signal ICO_DATA1_intermed_1 : std_logic_vector(31 downto 0);
signal R_M_CTRL_PC31DOWNTO12_intermed_4 : std_logic_vector(31 downto 12);
signal V_M_CTRL_TT3DOWNTO0_shadow_intermed_1 : std_logic_vector(3 downto 0);
signal V_X_CTRL_TT3DOWNTO0_shadow_intermed_1 : std_logic_vector(3 downto 0);
signal RIN_D_MEXC_intermed_3 : STD_ULOGIC;
signal V_E_CTRL_INST24_shadow_intermed_1 : STD_LOGIC;
signal R_W_S_TT3DOWNTO0_intermed_2 : STD_LOGIC_VECTOR(3 downto 0);
signal DSUIN_CRDY2_intermed_2 : STD_LOGIC;
signal V_X_RESULT6DOWNTO0_shadow_intermed_2 : std_logic_vector(6 downto 0);
signal RIN_D_PC3DOWNTO2_intermed_2 : std_logic_vector(3 downto 2);
signal V_D_PC_shadow_intermed_1 : std_logic_vector(31 downto 2);
signal R_A_CTRL_PC31DOWNTO4_intermed_2 : std_logic_vector(31 downto 4);
signal RIN_E_CTRL_RD6DOWNTO0_intermed_3 : std_logic_vector(6 downto 0);
signal R_A_CTRL_PC31DOWNTO12_intermed_4 : std_logic_vector(31 downto 12);
signal V_X_DATA031_shadow_intermed_1 : STD_LOGIC;
signal RIN_X_ANNUL_ALL_intermed_2 : STD_ULOGIC;
signal IRIN_ADDR3DOWNTO2_intermed_2 : std_logic_vector(3 downto 2);
signal RIN_D_SET_intermed_1 : STD_LOGIC_VECTOR(0 downto 0);
signal DCO_DATA0_intermed_1 : std_logic_vector(31 downto 0);
signal R_E_CTRL_CNT_intermed_2 : std_logic_vector(1 downto 0);
signal RIN_W_S_S_intermed_2 : STD_ULOGIC;
signal IRIN_ADDR31DOWNTO12_intermed_1 : std_logic_vector(31 downto 12);
signal RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_3 : std_logic_vector(3 downto 0);
signal RIN_W_S_TT3DOWNTO0_intermed_2 : STD_LOGIC_VECTOR(3 downto 0);
signal V_A_CTRL_LD_shadow_intermed_3 : STD_ULOGIC;
signal V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 : std_logic_vector(31 downto 2);
signal RIN_M_CTRL_PC_intermed_2 : std_logic_vector(31 downto 2);
signal R_D_INST1_intermed_2 : std_logic_vector(31 downto 0);
signal V_E_CTRL_shadow_intermed_2 : PIPELINE_CTRL_TYPE;
signal RIN_X_DATA1_intermed_1 : std_logic_vector(31 downto 0);
signal RIN_A_SU_intermed_2 : STD_ULOGIC;
signal R_A_CTRL_RD6DOWNTO0_intermed_2 : std_logic_vector(6 downto 0);
signal RIN_A_CTRL_PC31DOWNTO2_intermed_3 : std_logic_vector(31 downto 2);
signal RIN_E_CTRL_intermed_1 : PIPELINE_CTRL_TYPE;
signal RIN_A_CTRL_RD6DOWNTO0_intermed_3 : std_logic_vector(6 downto 0);
signal RIN_A_CTRL_TT3DOWNTO0_intermed_1 : std_logic_vector(3 downto 0);
signal RIN_F_PC_intermed_1 : std_logic_vector(31 downto 2);
signal V_D_PC31DOWNTO2_shadow_intermed_8 : std_logic_vector(31 downto 2);
signal V_D_CNT_shadow_intermed_1 : std_logic_vector(1 downto 0);
signal RIN_A_CTRL_LD_intermed_2 : STD_ULOGIC;
signal V_D_PC31DOWNTO4_shadow_intermed_5 : std_logic_vector(31 downto 4);
signal RIN_M_CTRL_PC31DOWNTO4_intermed_4 : std_logic_vector(31 downto 4);
signal R_A_CTRL_RETT_intermed_1 : STD_ULOGIC;
signal RIN_E_CTRL_INST_intermed_3 : std_logic_vector(31 downto 0);
signal R_D_MEXC_intermed_4 : STD_ULOGIC;
signal RIN_M_RESULT1DOWNTO0_intermed_3 : std_logic_vector(1 downto 0);
signal RIN_D_CNT_intermed_5 : std_logic_vector(1 downto 0);
signal V_A_CTRL_PC31DOWNTO12_shadow_intermed_1 : std_logic_vector(31 downto 12);
signal R_D_PC31DOWNTO2_intermed_3 : std_logic_vector(31 downto 2);
signal RIN_M_CTRL_PC31DOWNTO12_intermed_4 : std_logic_vector(31 downto 12);
signal RIN_M_CTRL_TT3DOWNTO0_intermed_1 : std_logic_vector(3 downto 0);
signal RIN_D_ANNUL_intermed_1 : STD_ULOGIC;
signal V_A_CTRL_shadow_intermed_1 : PIPELINE_CTRL_TYPE;
signal V_E_CTRL_PC31DOWNTO12_shadow_intermed_1 : std_logic_vector(31 downto 12);
signal RIN_M_CTRL_PC3DOWNTO2_intermed_4 : std_logic_vector(3 downto 2);
signal V_A_CTRL_PC31DOWNTO12_shadow_intermed_5 : std_logic_vector(31 downto 12);
signal R_D_PC31DOWNTO2_intermed_2 : std_logic_vector(31 downto 2);
signal RIN_E_CTRL_PC3DOWNTO2_intermed_5 : std_logic_vector(3 downto 2);
signal RIN_E_CTRL_PC31DOWNTO12_intermed_1 : std_logic_vector(31 downto 12);
signal R_A_CTRL_PC_intermed_4 : std_logic_vector(31 downto 2);
signal R_A_CTRL_ANNUL_intermed_4 : STD_ULOGIC;
signal V_X_RESULT_shadow_intermed_1 : std_logic_vector(31 downto 0);
signal R_E_CTRL_PC31DOWNTO2_intermed_1 : std_logic_vector(31 downto 2);
signal R_A_CTRL_PC31DOWNTO4_intermed_3 : std_logic_vector(31 downto 4);
signal V_D_CNT_shadow_intermed_5 : std_logic_vector(1 downto 0);
signal R_A_CTRL_TT_intermed_2 : std_logic_vector(5 downto 0);
signal RIN_A_CTRL_PC31DOWNTO12_intermed_5 : std_logic_vector(31 downto 12);
signal V_A_CTRL_TT3DOWNTO0_shadow_intermed_5 : std_logic_vector(3 downto 0);
signal RIN_W_S_S_intermed_1 : STD_ULOGIC;
signal V_M_CTRL_CNT_shadow_intermed_1 : std_logic_vector(1 downto 0);
signal V_A_CTRL_PC31DOWNTO12_shadow_intermed_7 : std_logic_vector(31 downto 12);
signal V_A_CTRL_WICC_shadow_intermed_2 : STD_ULOGIC;
signal R_X_DATA03_intermed_1 : STD_LOGIC;
signal RIN_M_DCI_intermed_1 : DC_IN_TYPE;
signal R_A_CTRL_CNT_intermed_2 : std_logic_vector(1 downto 0);
signal RIN_W_S_EF_intermed_1 : STD_ULOGIC;
signal V_E_CTRL_RD6DOWNTO0_shadow_intermed_2 : std_logic_vector(6 downto 0);
signal RIN_A_CTRL_LD_intermed_3 : STD_ULOGIC;
signal V_M_CTRL_RD6DOWNTO0_shadow_intermed_1 : std_logic_vector(6 downto 0);
signal R_E_CTRL_INST_intermed_2 : std_logic_vector(31 downto 0);
signal RIN_M_CTRL_RD6DOWNTO0_intermed_1 : std_logic_vector(6 downto 0);
signal V_F_PC3DOWNTO2_shadow_intermed_1 : std_logic_vector(3 downto 2);
signal EX_ADD_RES32DOWNTO330DOWNTO11_shadow_intermed_2 : STD_LOGIC_VECTOR(30 downto 11);
signal V_X_ANNUL_ALL_shadow_intermed_3 : STD_ULOGIC;
signal V_F_PC31DOWNTO12_shadow_intermed_2 : std_logic_vector(31 downto 12);
signal RIN_E_CTRL_INST24_intermed_1 : STD_LOGIC;
signal R_A_CTRL_PV_intermed_1 : STD_ULOGIC;
signal RIN_A_CTRL_RETT_intermed_3 : STD_ULOGIC;
signal R_E_CTRL_TT_intermed_2 : std_logic_vector(5 downto 0);
signal RIN_D_PC31DOWNTO12_intermed_7 : std_logic_vector(31 downto 12);
signal EX_ADD_RES32DOWNTO34DOWNTO3_shadow_intermed_1 : STD_LOGIC_VECTOR(4 downto 3);
signal V_E_CTRL_INST_shadow_intermed_2 : std_logic_vector(31 downto 0);
signal V_M_CTRL_PC31DOWNTO12_shadow_intermed_1 : std_logic_vector(31 downto 12);
signal DCO_MEXC_intermed_1 : STD_ULOGIC;
signal RIN_E_CWP_intermed_1 : std_logic_vector(2 downto 0);
signal V_A_CTRL_CNT_shadow_intermed_4 : std_logic_vector(1 downto 0);
signal V_A_CTRL_ANNUL_shadow_intermed_2 : STD_ULOGIC;
signal R_A_CTRL_PC31DOWNTO12_intermed_3 : std_logic_vector(31 downto 12);
signal R_A_CTRL_PC31DOWNTO2_intermed_4 : std_logic_vector(31 downto 2);
signal R_X_RESULT6DOWNTO0_intermed_2 : std_logic_vector(6 downto 0);
signal RIN_A_SU_intermed_1 : STD_ULOGIC;
signal R_E_CTRL_intermed_1 : PIPELINE_CTRL_TYPE;
signal V_E_OP231_shadow_intermed_1 : STD_LOGIC;
signal RIN_A_CTRL_WREG_intermed_3 : STD_ULOGIC;
signal V_A_CTRL_INST_shadow_intermed_4 : std_logic_vector(31 downto 0);
signal V_E_CTRL_PC31DOWNTO12_shadow_intermed_6 : std_logic_vector(31 downto 12);
signal V_M_CTRL_PC3DOWNTO2_shadow_intermed_1 : std_logic_vector(3 downto 2);
signal RPIN_ERROR_intermed_2 : STD_ULOGIC;
signal R_E_CTRL_TT3DOWNTO0_intermed_3 : std_logic_vector(3 downto 0);
signal V_D_CWP_shadow_intermed_1 : std_logic_vector(2 downto 0);
signal V_E_CTRL_PC31DOWNTO2_shadow_intermed_4 : std_logic_vector(31 downto 2);
signal RIN_A_CTRL_PV_intermed_3 : STD_ULOGIC;
signal RIN_M_CTRL_PC31DOWNTO4_intermed_1 : std_logic_vector(31 downto 4);
signal RIN_E_CTRL_INST24_intermed_2 : STD_LOGIC;
signal RIN_X_DCI_SIZE_intermed_1 : std_logic_vector(1 downto 0);
signal RIN_F_PC31DOWNTO12_intermed_1 : std_logic_vector(31 downto 12);
signal R_A_CTRL_TT3DOWNTO0_intermed_3 : std_logic_vector(3 downto 0);
signal DCO_DATA00_intermed_1 : STD_LOGIC;
signal V_M_Y31_shadow_intermed_1 : STD_LOGIC;
signal R_E_CTRL_PC31DOWNTO2_intermed_5 : std_logic_vector(31 downto 2);
signal R_A_CTRL_PC31DOWNTO2_intermed_1 : std_logic_vector(31 downto 2);
signal V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 : std_logic_vector(31 downto 2);
signal R_A_CTRL_INST19_intermed_1 : STD_LOGIC;
signal RIN_E_CTRL_TT_intermed_1 : std_logic_vector(5 downto 0);
signal RIN_E_CTRL_PC31DOWNTO2_intermed_2 : std_logic_vector(31 downto 2);
signal R_X_CTRL_PC3DOWNTO2_intermed_2 : std_logic_vector(3 downto 2);
signal RIN_X_ANNUL_ALL_intermed_4 : STD_ULOGIC;
signal V_A_CTRL_INST_shadow_intermed_1 : std_logic_vector(31 downto 0);
signal V_X_CTRL_PC31DOWNTO12_shadow_intermed_2 : std_logic_vector(31 downto 12);
signal IRIN_ADDR31DOWNTO4_intermed_2 : std_logic_vector(31 downto 4);
signal RIN_E_CTRL_PC3DOWNTO2_intermed_4 : std_logic_vector(3 downto 2);
signal RIN_A_CTRL_PC31DOWNTO4_intermed_1 : std_logic_vector(31 downto 4);
signal DCO_DATA04DOWNTO0_intermed_1 : std_logic_vector(4 downto 0);
signal RIN_E_CTRL_ANNUL_intermed_2 : STD_ULOGIC;
signal V_E_CTRL_INST19_shadow_intermed_1 : STD_LOGIC;
signal RIN_A_CTRL_PC_intermed_3 : std_logic_vector(31 downto 2);
signal V_X_DATA03_shadow_intermed_1 : STD_LOGIC;
signal V_E_OP1_shadow_intermed_1 : std_logic_vector(31 downto 0);
signal RIN_M_CTRL_CNT_intermed_2 : std_logic_vector(1 downto 0);
signal RIN_A_CTRL_PC31DOWNTO2_intermed_6 : std_logic_vector(31 downto 2);
signal RIN_D_MEXC_intermed_2 : STD_ULOGIC;
signal R_D_PC31DOWNTO4_intermed_2 : std_logic_vector(31 downto 4);
signal RIN_X_CTRL_INST_intermed_1 : std_logic_vector(31 downto 0);
signal V_A_SU_shadow_intermed_2 : STD_ULOGIC;
signal V_M_Y31_shadow_intermed_2 : STD_LOGIC;
signal R_W_S_TT3DOWNTO0_intermed_1 : STD_LOGIC_VECTOR(3 downto 0);
signal R_A_CTRL_ANNUL_intermed_3 : STD_ULOGIC;
signal R_A_CTRL_TRAP_intermed_1 : STD_ULOGIC;
signal RIN_M_CTRL_WICC_intermed_1 : STD_ULOGIC;
signal R_D_PC31DOWNTO2_intermed_7 : std_logic_vector(31 downto 2);
signal RIN_X_ANNUL_ALL_intermed_1 : STD_ULOGIC;
signal V_M_CTRL_WREG_shadow_intermed_1 : STD_ULOGIC;
signal V_A_CTRL_RD7DOWNTO0_shadow_intermed_4 : std_logic_vector(7 downto 0);
signal RIN_A_RFE1_intermed_1 : STD_ULOGIC;
signal V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 : std_logic_vector(31 downto 2);
signal V_D_PC31DOWNTO4_shadow_intermed_4 : std_logic_vector(31 downto 4);
signal R_A_CTRL_PC31DOWNTO12_intermed_2 : std_logic_vector(31 downto 12);
signal V_M_MAC_shadow_intermed_1 : STD_ULOGIC;
signal V_D_PC31DOWNTO2_shadow_intermed_2 : std_logic_vector(31 downto 2);
signal RIN_A_CTRL_TRAP_intermed_2 : STD_ULOGIC;
signal R_E_CTRL_RD7DOWNTO0_intermed_1 : std_logic_vector(7 downto 0);
signal R_E_CTRL_PC_intermed_3 : std_logic_vector(31 downto 2);
signal R_X_DATA00_intermed_1 : STD_LOGIC;
signal V_X_ANNUL_ALL_shadow_intermed_1 : STD_ULOGIC;
signal R_D_PC_intermed_5 : std_logic_vector(31 downto 2);
signal R_X_DATA03_intermed_2 : STD_LOGIC;
signal RIN_F_PC31DOWNTO4_intermed_1 : std_logic_vector(31 downto 4);
signal RIN_W_S_CWP_intermed_1 : std_logic_vector(2 downto 0);
signal V_W_S_PS_shadow_intermed_1 : STD_ULOGIC;
signal R_A_CTRL_intermed_1 : PIPELINE_CTRL_TYPE;
signal R_A_CTRL_TT_intermed_3 : std_logic_vector(5 downto 0);
signal RIN_A_CTRL_PC31DOWNTO4_intermed_6 : std_logic_vector(31 downto 4);
signal V_D_PC31DOWNTO2_shadow_intermed_7 : std_logic_vector(31 downto 2);
signal RIN_M_CTRL_PC31DOWNTO2_intermed_1 : std_logic_vector(31 downto 2);
signal R_X_DATA1_intermed_2 : std_logic_vector(31 downto 0);
signal R_D_PC3DOWNTO2_intermed_1 : std_logic_vector(3 downto 2);
signal RIN_X_CTRL_PC3DOWNTO2_intermed_1 : std_logic_vector(3 downto 2);
signal V_E_MAC_shadow_intermed_1 : STD_ULOGIC;
signal RIN_X_ICC_intermed_1 : STD_LOGIC_VECTOR(3 downto 0);
signal RIN_M_MAC_intermed_1 : STD_ULOGIC;
signal RIN_W_S_TT3DOWNTO0_intermed_1 : STD_LOGIC_VECTOR(3 downto 0);
signal R_D_PC31DOWNTO4_intermed_4 : std_logic_vector(31 downto 4);
signal V_A_CTRL_PC3DOWNTO2_shadow_intermed_6 : std_logic_vector(3 downto 2);
signal R_X_ANNUL_ALL_intermed_1 : STD_ULOGIC;
signal EX_JUMP_ADDRESS_shadow_intermed_1 : std_logic_vector(31 downto 2);
signal RIN_X_CTRL_PV_intermed_1 : STD_ULOGIC;
signal EX_ADD_RES32DOWNTO332DOWNTO13_shadow_intermed_2 : STD_LOGIC_VECTOR(32 downto 13);
signal RIN_A_CTRL_INST_intermed_1 : std_logic_vector(31 downto 0);
signal R_A_CTRL_RD6DOWNTO0_intermed_3 : std_logic_vector(6 downto 0);
signal IR_ADDR31DOWNTO12_intermed_1 : std_logic_vector(31 downto 12);
signal RIN_D_PC3DOWNTO2_intermed_6 : std_logic_vector(3 downto 2);
signal RIN_M_Y31_intermed_2 : STD_LOGIC;
signal RIN_X_DATA04DOWNTO0_intermed_2 : std_logic_vector(4 downto 0);
signal V_D_PC31DOWNTO2_shadow_intermed_3 : std_logic_vector(31 downto 2);
signal R_M_DCI_SIZE_intermed_1 : std_logic_vector(1 downto 0);
signal V_E_CTRL_PC3DOWNTO2_shadow_intermed_4 : std_logic_vector(3 downto 2);
signal V_E_OP2_shadow_intermed_1 : std_logic_vector(31 downto 0);
signal V_E_CTRL_TT3DOWNTO0_shadow_intermed_5 : std_logic_vector(3 downto 0);
signal V_A_CTRL_INST20_shadow_intermed_2 : STD_LOGIC;
signal RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1 : std_logic_vector(3 downto 0);
signal V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_4 : std_logic_vector(3 downto 0);
signal R_X_RESULT6DOWNTO03DOWNTO0_intermed_2 : std_logic_vector(3 downto 0);
signal RIN_M_CTRL_TRAP_intermed_2 : STD_ULOGIC;
signal V_A_CTRL_INST_shadow_intermed_3 : std_logic_vector(31 downto 0);


begin

  comb : process(ico, dco, rfo, r, wpr, ir, dsur, rstn, holdn, irqi, dbgi, fpo, cpo, tbo,
		 mulo, divo, dummy, rp)

  variable v 	: registers;
  variable vp 	: pwd_register_type;
  variable vwpr : watchpoint_registers;
  variable vdsu : dsu_registers;
  variable npc 	: std_logic_vector(31 downto 2);
  variable de_raddr1, de_raddr2 : std_logic_vector(9 downto 0);
  variable de_rs2, de_rd : std_logic_vector(4 downto 0);
  variable de_hold_pc, de_branch, de_fpop, de_ldlock : std_ulogic;
  variable de_cwp, de_cwp2 : cwptype;
  variable de_inull : std_ulogic;
  variable de_ren1, de_ren2 : std_ulogic;
  variable de_wcwp : std_ulogic;
  variable de_inst : word;
  variable de_branch_address : pctype;
  variable de_icc : std_logic_vector(3 downto 0);
  variable de_fbranch, de_cbranch : std_ulogic;
  variable de_rs1mod : std_ulogic;

  variable ra_op1, ra_op2 : word;
  variable ra_div : std_ulogic;

  variable ex_jump, ex_link_pc : std_ulogic;
  variable ex_jump_address : pctype;
  variable ex_add_res : std_logic_vector(32 downto 0);
  variable ex_shift_res, ex_logic_res, ex_misc_res : word;
  variable ex_edata, ex_edata2 : word;
  variable ex_dci : dc_in_type;
  variable ex_force_a2, ex_load, ex_ymsb : std_ulogic;
  variable ex_op1, ex_op2, ex_result, ex_result2, mul_op2 : word;
  variable ex_shcnt : std_logic_vector(4 downto 0);
  variable ex_dsuen : std_ulogic;
  variable ex_ldbp2 : std_ulogic;
  variable ex_sari : std_ulogic;
  
  variable me_inull, me_nullify, me_nullify2 : std_ulogic;
  variable me_iflush : std_ulogic;
  variable me_newtt : std_logic_vector(5 downto 0);
  variable me_asr18 : word;
  variable me_signed : std_ulogic;
  variable me_size, me_laddr : std_logic_vector(1 downto 0);
  variable me_icc : std_logic_vector(3 downto 0);

  
  variable xc_result : word;
  variable xc_df_result : word;
  variable xc_waddr : std_logic_vector(9 downto 0);
  variable xc_exception, xc_wreg : std_ulogic;
  variable xc_trap_address : pctype;
  variable xc_vectt : std_logic_vector(7 downto 0);
  variable xc_trap : std_ulogic;
  variable xc_fpexack : std_ulogic;
  variable xc_rstn, xc_halt : std_ulogic;
  
--  variable wr_rf1_data, wr_rf2_data : word;
  variable diagdata : word;
  variable tbufi : tracebuf_in_type;
  variable dbgm : std_ulogic;
  variable fpcdbgwr : std_ulogic;
  variable vfpi : fpc_in_type;
  variable dsign : std_ulogic;
  variable pwrd, sidle : std_ulogic;
  variable vir : irestart_register;
  variable icnt : std_ulogic;
  variable tbufcntx : std_logic_vector(7-1 downto 0);
  
  begin

    v := r; vwpr := wpr; vdsu := dsur; vp := rp;
    xc_fpexack := '0'; sidle := '0';
    fpcdbgwr := '0'; vir := ir; xc_rstn := rstn;
    
-----------------------------------------------------------------------
-- WRITE STAGE
-----------------------------------------------------------------------

--    wr_rf1_data := rfo.data1; wr_rf2_data := rfo.data2;
--    if irfwt = 0 then
--      if r.w.wreg = '1' then
--	if r.a.rfa1 = r.w.wa then wr_rf1_data := r.w.result; end if;
--	if r.a.rfa2 = r.w.wa then wr_rf2_data := r.w.result; end if;
--      end if;
--    end if;

-----------------------------------------------------------------------
-- EXCEPTION STAGE
-----------------------------------------------------------------------

    xc_exception := '0'; xc_halt := '0'; icnt := '0';
    xc_waddr := "0000000000";
    xc_waddr(7 downto 0) := r.x.ctrl.rd(7 downto 0);
    xc_trap := r.x.mexc or r.x.ctrl.trap;
    v.x.nerror := rp.error;
    
    if r.x.mexc = '1' then
      xc_vectt := "00" & TT_DAEX;
    elsif r.x.ctrl.tt = TT_TICC then
      xc_vectt := '1' & r.x.result(6 downto 0);
    else xc_vectt := "00" & r.x.ctrl.tt; end if;
    if r.w.s.svt = '0' then
      xc_trap_address(31 downto 4) := r.w.s.tba & xc_vectt; 
    else
      xc_trap_address(31 downto 4) := r.w.s.tba & "00000000"; 
    end if;
    xc_trap_address(3 downto 2) := "00";
    xc_wreg := '0'; v.x.annul_all := '0'; 
    if (r.x.ctrl.ld = '1') then 
      if (lddel = 2) then 
        xc_result := ld_align(r.x.data, r.x.set, r.x.dci.size, r.x.laddr, r.x.dci.signed);
      else xc_result := r.x.data(0); end if;
    elsif false and false and (r.x.mac = '1') then
      xc_result := mulo.result(31 downto 0);
    else xc_result := r.x.result; end if;
    xc_df_result := xc_result;
    if true then 
      dbgm := dbgexc(r, dbgi, xc_trap, xc_vectt);
      if (dbgi.dsuen and dbgi.dbreak) = '0'then v.x.debug := '0'; end if;
    else dbgm := '0'; v.x.debug := '0'; end if;
    if false then pwrd := powerdwn(r, xc_trap, rp); else pwrd := '0'; end if;
    
    case r.x.rstate is
    when run =>
      if (not r.x.ctrl.annul and r.x.ctrl.pv and not r.x.debug) = '1' then
	icnt := holdn;
      end if;
      if dbgm = '1' then        
        v.x.annul_all := '1'; vir.addr := r.x.ctrl.pc;
        v.x.rstate := dsu1; v.x.debug := '1';
        v.x.npc := npc_find(r);
        vdsu.tt := xc_vectt; vdsu.err := dbgerr(r, dbgi, xc_vectt);
      elsif (pwrd = '1') and (ir.pwd = '0') then
        v.x.annul_all := '1'; vir.addr := r.x.ctrl.pc;
        v.x.rstate := dsu1; v.x.npc := npc_find(r); vp.pwd := '1';
      elsif (r.x.ctrl.annul or xc_trap) = '0' then
        xc_wreg := r.x.ctrl.wreg;
        sp_write (r, wpr, v.w.s, vwpr);        
        vir.pwd := '0';
      elsif ((not r.x.ctrl.annul) and xc_trap) = '1' then
        xc_exception := '1'; xc_result := r.x.ctrl.pc(31 downto 2) & "00";
        xc_wreg := '1'; v.w.s.tt := xc_vectt; v.w.s.ps := r.w.s.s;
        v.w.s.s := '1'; v.x.annul_all := '1'; v.x.rstate := trap;
        xc_waddr := "0000000000";
        xc_waddr(6  downto 0) :=  r.w.s.cwp & "0001";
	v.x.npc := npc_find(r);
        fpexack(r, xc_fpexack);
        if r.w.s.et = '0' then
--	  v.x.rstate := dsu1; xc_wreg := '0'; vp.error := '1';
	   xc_wreg := '0';
        end if;
      end if;
    when trap =>
      xc_result := npc_gen(r); xc_wreg := '1';
      xc_waddr := "0000000000";
      xc_waddr(6  downto 0) :=  r.w.s.cwp & "0010";
      if (r.w.s.et = '1') then
	v.w.s.et := '0'; v.x.rstate := run;
        if (not true) and (r.w.s.cwp = "000") then v.w.s.cwp := "111";
        else v.w.s.cwp := r.w.s.cwp - 1 ; end if;
      else
	v.x.rstate := dsu1; xc_wreg := '0'; vp.error := '1';
      end if;
    when dsu1 =>
      xc_exception := '1'; v.x.annul_all := '1';
      xc_trap_address(31 downto 2) := r.f.pc;        
      if true or false or (smp /= 0) then 
        xc_trap_address(31 downto 2) := ir.addr; 
        vir.addr := npc_gen(r)(31 downto 2);
        v.x.rstate := dsu2;
      end if;
      if true then v.x.debug := r.x.debug; end if;
    when dsu2 =>      
      xc_exception := '1'; v.x.annul_all := '1';
      xc_trap_address(31 downto 2) := r.f.pc;        
      if true or false or (smp /= 0) then
	sidle := (rp.pwd or rp.error) and ico.idle and dco.idle and not r.x.debug;
        if true then
	  if dbgi.reset = '1' then 
	    if smp /=0 then vp.pwd := not irqi.run; else vp.pwd := '0'; end if;
	    vp.error := '0';
	  end if;
          if (dbgi.dsuen and dbgi.dbreak) = '1'then v.x.debug := '1'; end if;
          diagwr(r, dsur, ir, dbgi, wpr, v.w.s, vwpr, vdsu.asi, xc_trap_address,
            vir.addr, vdsu.tbufcnt, xc_wreg, xc_waddr, xc_result, fpcdbgwr);
	  xc_halt := dbgi.halt;
        end if;
	if r.x.ipend = '1' then vp.pwd := '0'; end if;
        if (rp.error or rp.pwd or r.x.debug or xc_halt) = '0' then
	  v.x.rstate := run; v.x.annul_all := '0'; vp.error := '0';
          xc_trap_address(31 downto 2) := ir.addr; v.x.debug := '0';
          vir.pwd := '1';
        end if;
        if (smp /= 0) and (irqi.rst = '1') then 
	  vp.pwd := '0'; vp.error := '0';
	end if;
      end if;
    when others =>
    end case;

    irq_intack(r, holdn, v.x.intack);          
    itrace(r, dsur, vdsu, xc_result, xc_exception, dbgi, rp.error, xc_trap, tbufcntx, tbufi);
    vdsu.tbufcnt := tbufcntx;

    v.w.except := xc_exception; v.w.result := xc_result;
    if (r.x.rstate = dsu2) then v.w.except := '0'; end if;
    v.w.wa := xc_waddr(7 downto 0); v.w.wreg := xc_wreg and holdn;

    rfi.wdata <= xc_result; rfi.waddr <= xc_waddr;
    rfi.wren <= (xc_wreg and holdn) and not dco.scanen;
    irqo.intack <= r.x.intack and holdn;
    irqo.irl <= r.w.s.tt(3 downto 0);
    irqo.pwd <= rp.pwd;
    irqo.fpen <= r.w.s.ef;
    dbgo.halt <= xc_halt;
    dbgo.pwd <= rp.pwd;
    dbgo.idle <= sidle;
    dbgo.icnt <= icnt;
    dci.intack <= r.x.intack and holdn;
    
    if (xc_rstn = '0') then 
      v.w.except := '0'; v.w.s.et := '0'; v.w.s.svt := '0'; v.w.s.dwt := '0';
      v.w.s.ef := '0';  -- needed for AX
      if need_extra_sync_reset(fabtech) /= 0 then 
	v.w.s.cwp := "000";
	v.w.s.icc := "0000";
      end if;
      v.x.annul_all := '1'; v.x.rstate := run; vir.pwd := '0'; 
      vp.pwd := '0'; v.x.debug := '0'; --vp.error := '0';
      v.x.nerror := '0';
      if svt = 1 then  v.w.s.tt := "00000000"; end if;
      if true then
        if (dbgi.dsuen and dbgi.dbreak) = '1' then
          v.x.rstate := dsu1; v.x.debug := '1';
        end if;
      end if;
      if (smp /= 0) and (irqi.run = '0') and (rstn = '0') then 
	v.x.rstate := dsu1; vp.pwd := '1';
      end if;
    end if;
    
    if not FPEN then v.w.s.ef := '0'; end if;

-----------------------------------------------------------------------
-- MEMORY STAGE
-----------------------------------------------------------------------

    v.x.ctrl := r.m.ctrl; v.x.dci := r.m.dci;
    v.x.ctrl.rett := r.m.ctrl.rett and not r.m.ctrl.annul;
    v.x.mac := r.m.mac; v.x.laddr := r.m.result(1 downto 0);
    v.x.ctrl.annul := r.m.ctrl.annul or v.x.annul_all; 
    
    mul_res(r, v.w.s.asr18, v.x.result, v.x.y, me_asr18, me_icc);
    mem_trap(r, wpr, v.x.ctrl.annul, holdn, v.x.ctrl.trap, me_iflush,
	     me_nullify, v.m.werr, v.x.ctrl.tt);
    me_newtt := v.x.ctrl.tt;

    irq_trap(r, ir, irqi.irl, v.x.ctrl.annul, v.x.ctrl.pv, v.x.ctrl.trap, me_newtt, me_nullify,
             v.m.irqen, v.m.irqen2, me_nullify2, v.x.ctrl.trap,
	     v.x.ipend, v.x.ctrl.tt);   
    
    if (r.m.ctrl.ld or not dco.mds) = '1' then 
      for i in 0 to 2-1 loop v.x.data(i) := dco.data(i); end loop;
      v.x.set := dco.set(0 downto 0);
      if dco.mds = '0' then
	me_size := r.x.dci.size; me_laddr := r.x.laddr; me_signed := r.x.dci.signed;
      else
	me_size := v.x.dci.size; me_laddr := v.x.laddr; me_signed := v.x.dci.signed;
      end if;
      if lddel /= 2 then
        v.x.data(0) := ld_align(v.x.data, v.x.set, me_size, me_laddr, me_signed);
      end if;
    end if;
    v.x.mexc := dco.mexc;

    v.x.icc := me_icc;
    v.x.ctrl.wicc := r.m.ctrl.wicc and not v.x.annul_all;
    
    if false and ((v.x.ctrl.annul or v.x.ctrl.trap) = '0') then
      v.w.s.asr18 := me_asr18;
    end if;

    if (r.x.rstate = dsu2) then
      me_nullify2 := '0'; v.x.set := dco.set(0 downto 0);
    end if;

    dci.maddress <= r.m.result;
    dci.msu    <= r.m.su;
    dci.esu    <= r.e.su;
    dci.enaddr   <= r.m.dci.enaddr;
    dci.asi      <= r.m.dci.asi;
    dci.size     <= r.m.dci.size;
    dci.nullify  <= me_nullify2;
    dci.lock     <= r.m.dci.lock and not r.m.ctrl.annul;
    dci.read     <= r.m.dci.read;
    dci.write    <= r.m.dci.write;
    dci.flush    <= me_iflush;
    dci.dsuen    <= r.m.dci.dsuen;
    dbgo.ipend <= v.x.ipend;

-----------------------------------------------------------------------
-- EXECUTE STAGE
-----------------------------------------------------------------------

    v.m.ctrl := r.e.ctrl; ex_op1 := r.e.op1; ex_op2 := r.e.op2;
    v.m.ctrl.rett := r.e.ctrl.rett and not r.e.ctrl.annul;
    v.m.ctrl.wreg := r.e.ctrl.wreg and not v.x.annul_all;    
    ex_ymsb := r.e.ymsb; mul_op2 := ex_op2; ex_shcnt := r.e.shcnt;
    v.e.cwp := r.a.cwp; ex_sari := r.e.sari;
    v.m.su := r.e.su;
    if 0 = 3 then v.m.mul := r.e.mul; else v.m.mul := '0'; end if;

    if lddel = 1 then
      if r.e.ldbp1 = '1' then 
	ex_op1 := r.x.data(0); 
	ex_sari := r.x.data(0)(31) and r.e.ctrl.inst(19) and r.e.ctrl.inst(20);
      end if;
      if r.e.ldbp2 = '1' then 
	ex_op2 := r.x.data(0); ex_ymsb := r.x.data(0)(0); 
	mul_op2 := ex_op2; ex_shcnt := r.x.data(0)(4 downto 0);
	if r.e.invop2 = '1' then 
	  ex_op2 := not ex_op2; ex_shcnt := not ex_shcnt;
        end if;
      end if;
    end if;

    ex_add_res := (ex_op1 & '1') + (ex_op2 & r.e.alucin);

    if ex_add_res(2 downto 1) = "00" then v.m.nalign := '0';
    else v.m.nalign := '1'; end if;

    dcache_gen(r, v, ex_dci, ex_link_pc, ex_jump, ex_force_a2, ex_load );
    ex_jump_address := ex_add_res(32 downto 3);
    logic_op(r, ex_op1, ex_op2, v.x.y, ex_ymsb, ex_logic_res, v.m.y);
    ex_shift_res := shift(r, ex_op1, ex_op2, ex_shcnt, ex_sari);
    misc_op(r, wpr, ex_op1, ex_op2, xc_df_result, v.x.y, ex_misc_res, ex_edata);
    ex_add_res(3):= ex_add_res(3) or ex_force_a2;    
    alu_select(r, ex_add_res, ex_op1, ex_op2, ex_shift_res, ex_logic_res,
	ex_misc_res, ex_result, me_icc, v.m.icc, v.m.divz);    
    dbg_cache(holdn, dbgi, r, dsur, ex_result, ex_dci, ex_result2, v.m.dci);
    fpstdata(r, ex_edata, ex_result2, fpo.data, ex_edata2, v.m.result);
    cwp_ex(r, v.m.wcwp);    
    
    v.m.ctrl.annul := v.m.ctrl.annul or v.x.annul_all;
    v.m.ctrl.wicc := r.e.ctrl.wicc and not v.x.annul_all; 
    v.m.mac := r.e.mac;
    if (true and (r.x.rstate = dsu2)) then v.m.ctrl.ld := '1'; end if;
    dci.eenaddr  <= v.m.dci.enaddr;
    dci.eaddress <= ex_add_res(32 downto 1);
    dci.edata <= ex_edata2;
    
-----------------------------------------------------------------------
-- REGFILE STAGE
-----------------------------------------------------------------------

    v.e.ctrl := r.a.ctrl; v.e.jmpl := r.a.jmpl;
    v.e.ctrl.annul := r.a.ctrl.annul or v.x.annul_all;
    v.e.ctrl.rett := r.a.ctrl.rett and not r.a.ctrl.annul;
    v.e.ctrl.wreg := r.a.ctrl.wreg and not v.x.annul_all;    
    v.e.su := r.a.su; v.e.et := r.a.et;
    v.e.ctrl.wicc := r.a.ctrl.wicc and not v.x.annul_all;
    
    exception_detect(r, wpr, dbgi, r.a.ctrl.trap, r.a.ctrl.tt, 
		     v.e.ctrl.trap, v.e.ctrl.tt);
    op_mux(r, rfo.data1, v.m.result, v.x.result, xc_df_result, "00000000000000000000000000000000", 
	r.a.rsel1, v.e.ldbp1, ra_op1);
    op_mux(r, rfo.data2,  v.m.result, v.x.result, xc_df_result, r.a.imm, 
	r.a.rsel2, ex_ldbp2, ra_op2);
    alu_op(r, ra_op1, ra_op2, v.m.icc, v.m.y(0), ex_ldbp2, v.e.op1, v.e.op2,
	   v.e.aluop, v.e.alusel, v.e.aluadd, v.e.shcnt, v.e.sari, v.e.shleft,
	   v.e.ymsb, v.e.mul, ra_div, v.e.mulstep, v.e.mac, v.e.ldbp2, v.e.invop2);
    cin_gen(r, v.m.icc(0), v.e.alucin);

-----------------------------------------------------------------------
-- DECODE STAGE
-----------------------------------------------------------------------

    if 2 > 1 then de_inst := r.d.inst(conv_integer(r.d.set));
    else de_inst := r.d.inst(0); end if;

    de_icc := r.m.icc; v.a.cwp := r.d.cwp;
    su_et_select(r, v.w.s.ps, v.w.s.s, v.w.s.et, v.a.su, v.a.et);
    wicc_y_gen(de_inst, v.a.ctrl.wicc, v.a.ctrl.wy);
    cwp_ctrl(r, v.w.s.wim, de_inst, de_cwp, v.a.wovf, v.a.wunf, de_wcwp);
    rs1_gen(r, de_inst, v.a.rs1, de_rs1mod); 
    de_rs2 := de_inst(4 downto 0);
    de_raddr1 := "0000000000"; de_raddr2 := "0000000000";
    
    if true then
      if de_rs1mod = '1' then
        regaddr(r.d.cwp, de_inst(29 downto 26) & v.a.rs1(0), de_raddr1(7 downto 0));
      else
        regaddr(r.d.cwp, de_inst(18 downto 15) & v.a.rs1(0), de_raddr1(7 downto 0));
      end if;
    else
      regaddr(r.d.cwp, v.a.rs1, de_raddr1(7 downto 0));
    end if;
    regaddr(r.d.cwp, de_rs2, de_raddr2(7 downto 0));
    v.a.rfa1 := de_raddr1(7 downto 0); 
    v.a.rfa2 := de_raddr2(7 downto 0); 

    rd_gen(r, de_inst, v.a.ctrl.wreg, v.a.ctrl.ld, de_rd);
    regaddr(de_cwp, de_rd, v.a.ctrl.rd);
    
    fpbranch(de_inst, fpo.cc, de_fbranch);
    fpbranch(de_inst, cpo.cc, de_cbranch);
    v.a.imm := imm_data(r, de_inst);
    lock_gen(r, de_rs2, de_rd, v.a.rfa1, v.a.rfa2, v.a.ctrl.rd, de_inst, 
	fpo.ldlock, v.e.mul, ra_div, v.a.ldcheck1, v.a.ldcheck2, de_ldlock, 
	v.a.ldchkra, v.a.ldchkex);
    ic_ctrl(r, de_inst, v.x.annul_all, de_ldlock, branch_true(de_icc, de_inst), 
	de_fbranch, de_cbranch, fpo.ccv, cpo.ccv, v.d.cnt, v.d.pc, de_branch,
	v.a.ctrl.annul, v.d.annul, v.a.jmpl, de_inull, v.d.pv, v.a.ctrl.pv,
	de_hold_pc, v.a.ticc, v.a.ctrl.rett, v.a.mulstart, v.a.divstart);

    cwp_gen(r, v, v.a.ctrl.annul, de_wcwp, de_cwp, v.d.cwp);    
    
    v.d.inull := ra_inull_gen(r, v);

    op_find(r, v.a.ldchkra, v.a.ldchkex, v.a.rs1, v.a.rfa1, 
	    false, v.a.rfe1, v.a.rsel1, v.a.ldcheck1);
    op_find(r, v.a.ldchkra, v.a.ldchkex, de_rs2, v.a.rfa2, 
	    imm_select(de_inst), v.a.rfe2, v.a.rsel2, v.a.ldcheck2);

    de_branch_address := branch_address(de_inst, r.d.pc);

    v.a.ctrl.annul := v.a.ctrl.annul or v.x.annul_all;    
    v.a.ctrl.wicc := v.a.ctrl.wicc and not v.a.ctrl.annul;
    v.a.ctrl.wreg := v.a.ctrl.wreg and not v.a.ctrl.annul;
    v.a.ctrl.rett := v.a.ctrl.rett and not v.a.ctrl.annul;
    v.a.ctrl.wy := v.a.ctrl.wy and not v.a.ctrl.annul;

    v.a.ctrl.trap := r.d.mexc;
    v.a.ctrl.tt := "000000";
    v.a.ctrl.inst := de_inst;
    v.a.ctrl.pc := r.d.pc;
    v.a.ctrl.cnt := r.d.cnt;
    v.a.step := r.d.step;

    if holdn = '0' then 
      de_raddr1(7 downto 0) := r.a.rfa1;
      de_raddr2(7 downto 0) := r.a.rfa2;
      de_ren1 := r.a.rfe1; de_ren2 := r.a.rfe2;
    else
      de_ren1 := v.a.rfe1; de_ren2 := v.a.rfe2;
    end if;

    if true then
      if ((dbgi.denable and not dbgi.dwrite) = '1') and (r.x.rstate = dsu2) then        
        de_raddr1(7 downto 0) := dbgi.daddr(9 downto 2); de_ren1 := '1';
      end if;
      v.d.step := dbgi.step and not r.d.annul;      
    end if;

    rfi.raddr1 <= de_raddr1; rfi.raddr2 <= de_raddr2;
    rfi.ren1 <= de_ren1 and not dco.scanen;
    rfi.ren2 <= de_ren2 and not dco.scanen;
    rfi.diag <= dco.testen & "000";
    ici.inull <= de_inull;
    ici.flush <= me_iflush;
    if (xc_rstn = '0') then
      v.d.cnt := "00";
      if need_extra_sync_reset(fabtech) /= 0 then 
	v.d.cwp := "000";
      end if;
    end if;


-----------------------------------------------------------------------
-- FETCH STAGE
-----------------------------------------------------------------------

    npc := r.f.pc;
    if (xc_rstn = '0') then
      v.f.pc := "000000000000000000000000000000"; v.f.branch := '0';
      if false then v.f.pc(31 downto 12) := irqi.rstvec;
      else
        v.f.pc(31 downto 12) := conv_std_logic_vector(rstaddr, 20);
      end if;
    elsif xc_exception = '1' then	-- exception
      v.f.branch := '1'; v.f.pc := xc_trap_address;
      npc := v.f.pc;
--    elsif (not ra_inull and de_hold_pc) = '1' then
    elsif de_hold_pc = '1' then
      v.f.pc := r.f.pc; v.f.branch := r.f.branch;
      if ex_jump = '1' then
        v.f.pc := ex_jump_address; v.f.branch := '1';
        npc := v.f.pc;
      end if;
    elsif ex_jump = '1' then
      v.f.pc := ex_jump_address; v.f.branch := '1';
      npc := v.f.pc;
    elsif de_branch = '1' then
      v.f.pc := branch_address(de_inst, r.d.pc); v.f.branch := '1';
      npc := v.f.pc;
    else
      v.f.branch := '0';
      v.f.pc(31 downto 2) := r.f.pc(31 downto 2) + 1;    -- Address incrementer
      npc := v.f.pc;
    end if;

    ici.dpc <= r.d.pc(31 downto 2) & "00";
    ici.fpc <= r.f.pc(31 downto 2) & "00";
    ici.rpc <= npc(31 downto 2) & "00";
    ici.fbranch <= r.f.branch;
    ici.rbranch <= v.f.branch;
    ici.su <= v.a.su;
    ici.fline <= "00000000000000000000000000000";
    ici.flushl <= '0';

    if (ico.mds and de_hold_pc) = '0' then 
      for i in 0 to 2-1 loop
        v.d.inst(i) := ico.data(i);			-- latch instruction
      end loop;
      v.d.set := ico.set(0 downto 0);             -- latch instruction
      v.d.mexc := ico.mexc;				-- latch instruction
    end if;

-----------------------------------------------------------------------
-----------------------------------------------------------------------

    if true then -- DSU diagnostic read    
      diagread(dbgi, r, dsur, ir, wpr, dco, tbo, diagdata);
      diagrdy(dbgi.denable, dsur, r.m.dci, dco.mds, ico, vdsu.crdy);
    end if;
    
-----------------------------------------------------------------------
-- OUTPUTS
-----------------------------------------------------------------------

    rin <= v; wprin <= vwpr; dsuin <= vdsu; irin <= vir;
    muli.start <= r.a.mulstart and not r.a.ctrl.annul;
    muli.signed <= r.e.ctrl.inst(19);
    muli.op1 <= (ex_op1(31) and r.e.ctrl.inst(19)) & ex_op1;
    muli.op2 <= (mul_op2(31) and r.e.ctrl.inst(19)) & mul_op2;
    muli.mac <= r.e.ctrl.inst(24);
    if false then muli.acc(39 downto 32) <= r.w.s.y(7 downto 0);
    else muli.acc(39 downto 32) <= r.x.y(7 downto 0); end if;
    muli.acc(31 downto 0) <= r.w.s.asr18;
    muli.flush <= r.x.annul_all;
    divi.start <= r.a.divstart and not r.a.ctrl.annul;
    divi.signed <= r.e.ctrl.inst(19);
    divi.flush <= r.x.annul_all;
    divi.op1 <= (ex_op1(31) and r.e.ctrl.inst(19)) & ex_op1;
    divi.op2 <= (ex_op2(31) and r.e.ctrl.inst(19)) & ex_op2;
    if (r.a.divstart and not r.a.ctrl.annul) = '1' then 
      dsign :=  r.a.ctrl.inst(19);
    else dsign := r.e.ctrl.inst(19); end if;
    divi.y <= (r.m.y(31) and dsign) & r.m.y;
    rpin <= vp;

    if true then
      dbgo.dsu <= '1'; dbgo.dsumode <= r.x.debug; dbgo.crdy <= dsur.crdy(2);
      dbgo.data <= diagdata;
      if true then tbi <= tbufi; else
        tbi.addr <= (others => '0'); tbi.data <= (others => '0');
        tbi.enable <= '0'; tbi.write <= (others => '0'); tbi.diag <= "0000";
      end if;
    else
      dbgo.dsu <= '0'; dbgo.data <= (others => '0'); dbgo.crdy  <= '0';
      dbgo.dsumode <= '0';
      tbi.addr <= (others => '0'); tbi.data <= (others => '0');
      tbi.enable <= '0'; tbi.write <= (others => '0'); tbi.diag <= "0000";
    end if;
    dbgo.error <= dummy and not r.x.nerror;

-- pragma translate_off
    if FPEN then
-- pragma translate_on
      vfpi.flush := v.x.annul_all; vfpi.exack := xc_fpexack; vfpi.a_rs1 := r.a.rs1; vfpi.d.inst := de_inst;
      vfpi.d.cnt := r.d.cnt; vfpi.d.annul := v.x.annul_all or r.d.annul; vfpi.d.trap := r.d.mexc;
      vfpi.d.pc(1 downto 0) := (others => '0'); vfpi.d.pc(31 downto 2) := r.d.pc(31 downto 2); 
      vfpi.d.pv := r.d.pv;
      vfpi.a.pc(1 downto 0) := (others => '0'); vfpi.a.pc(31 downto 2) := r.a.ctrl.pc(31 downto 2); 
      vfpi.a.inst := r.a.ctrl.inst; vfpi.a.cnt := r.a.ctrl.cnt; vfpi.a.trap := r.a.ctrl.trap;
      vfpi.a.annul := r.a.ctrl.annul; vfpi.a.pv := r.a.ctrl.pv;
      vfpi.e.pc(1 downto 0) := (others => '0'); vfpi.e.pc(31 downto 2) := r.e.ctrl.pc(31 downto 2); 
      vfpi.e.inst := r.e.ctrl.inst; vfpi.e.cnt := r.e.ctrl.cnt; vfpi.e.trap := r.e.ctrl.trap; vfpi.e.annul := r.e.ctrl.annul;
      vfpi.e.pv := r.e.ctrl.pv;
      vfpi.m.pc(1 downto 0) := (others => '0'); vfpi.m.pc(31 downto 2) := r.m.ctrl.pc(31 downto 2); 
      vfpi.m.inst := r.m.ctrl.inst; vfpi.m.cnt := r.m.ctrl.cnt; vfpi.m.trap := r.m.ctrl.trap; vfpi.m.annul := r.m.ctrl.annul;
      vfpi.m.pv := r.m.ctrl.pv;
      vfpi.x.pc(1 downto 0) := (others => '0'); vfpi.x.pc(31 downto 2) := r.x.ctrl.pc(31 downto 2); 
      vfpi.x.inst := r.x.ctrl.inst; vfpi.x.cnt := r.x.ctrl.cnt; vfpi.x.trap := xc_trap;
      vfpi.x.annul := r.x.ctrl.annul; vfpi.x.pv := r.x.ctrl.pv; vfpi.lddata := xc_df_result;--xc_result;
      if r.x.rstate = dsu2 then vfpi.dbg.enable := dbgi.denable;
      else vfpi.dbg.enable := '0'; end if;      
      vfpi.dbg.write := fpcdbgwr;
      vfpi.dbg.fsr := dbgi.daddr(22); -- IU reg access
      vfpi.dbg.addr := dbgi.daddr(6 downto 2);
      vfpi.dbg.data := dbgi.ddata;
      fpi <= vfpi;
      cpi <= vfpi;  -- dummy, just to kill some warnings ...
-- pragma translate_off
    end if;
-- pragma translate_on
-- Assignments to be moved with variables

-- These assignments must be moved to process COMB/
V_A_ET_shadow <= V.A.ET;
EX_ADD_RES32DOWNTO34DOWNTO3_shadow <= EX_ADD_RES ( 32 DOWNTO 3 )( 4 DOWNTO 3 );
ICNT_shadow <= ICNT;
EX_OP1_shadow <= EX_OP1;
V_M_CTRL_PC_shadow <= V.M.CTRL.PC;
V_E_CTRL_PC3DOWNTO2_shadow <= V.E.CTRL.PC( 3 DOWNTO 2 );
DE_REN1_shadow <= DE_REN1;
DE_INST_shadow <= DE_INST;
V_A_CTRL_CNT_shadow <= V.A.CTRL.CNT;
V_F_PC3DOWNTO2_shadow <= V.F.PC( 3 DOWNTO 2 );
V_W_S_TT_shadow <= V.W.S.TT;
V_X_RESULT6DOWNTO0_shadow <= V.X.RESULT ( 6 DOWNTO 0 );
EX_JUMP_ADDRESS3DOWNTO2_shadow <= EX_JUMP_ADDRESS( 3 DOWNTO 2 );
V_E_ALUCIN_shadow <= V.E.ALUCIN;
V_D_PC3DOWNTO2_shadow <= V.D.PC( 3 DOWNTO 2 );
V_A_CTRL_PV_shadow <= V.A.CTRL.PV;
V_E_CTRL_shadow <= V.E.CTRL;
V_M_CTRL_shadow <= V.M.CTRL;
V_M_RESULT1DOWNTO0_shadow <= V.M.RESULT ( 1 DOWNTO 0 );
EX_SHCNT_shadow <= EX_SHCNT;
V_M_DCI_SIZE_shadow <= V.M.DCI.SIZE;
V_X_CTRL_ANNUL_shadow <= V.X.CTRL.ANNUL;
V_X_MEXC_shadow <= V.X.MEXC;
TBUFCNTX_shadow <= TBUFCNTX;
V_A_CTRL_WY_shadow <= V.A.CTRL.WY;
NPC_shadow <= NPC;
V_M_CTRL_TT3DOWNTO0_shadow <= V.M.CTRL.TT( 3 DOWNTO 0 );
V_A_MULSTART_shadow <= V.A.MULSTART;
XC_VECTT3DOWNTO0_shadow <= XC_VECTT( 3 DOWNTO 0 );
V_E_CTRL_TT_shadow <= V.E.CTRL.TT;
DSIGN_shadow <= DSIGN;
V_E_CTRL_ANNUL_shadow <= V.E.CTRL.ANNUL;
EX_JUMP_ADDRESS_shadow <= EX_JUMP_ADDRESS;
V_A_CTRL_PC31DOWNTO12_shadow <= V.A.CTRL.PC( 31 DOWNTO 12 );
V_A_RFE1_shadow <= V.A.RFE1;
V_W_WA_shadow <= V.W.WA;
V_X_ANNUL_ALL_shadow <= V.X.ANNUL_ALL;
EX_YMSB_shadow <= EX_YMSB;
EX_ADD_RES_shadow <= EX_ADD_RES;
VIR_ADDR_shadow <= VIR.ADDR;
EX_JUMP_ADDRESS31DOWNTO12_shadow <= EX_JUMP_ADDRESS( 31 DOWNTO 12 );
V_W_S_CWP_shadow <= V.W.S.CWP;
V_D_INST0_shadow <= V.D.INST ( 0 );
V_A_CTRL_ANNUL_shadow <= V.A.CTRL.ANNUL;
V_X_DATA1_shadow <= V.X.DATA ( 1 );
VP_PWD_shadow <= VP.PWD;
V_M_CTRL_RD6DOWNTO0_shadow <= V.M.CTRL.RD( 6 DOWNTO 0 );
V_X_DATA00_shadow <= V.X.DATA ( 0 )( 0 );
V_M_CTRL_RETT_shadow <= V.M.CTRL.RETT;
V_X_CTRL_RETT_shadow <= V.X.CTRL.RETT;
V_X_CTRL_PC31DOWNTO12_shadow <= V.X.CTRL.PC( 31 DOWNTO 12 );
V_W_S_PS_shadow <= V.W.S.PS;
V_X_CTRL_TT_shadow <= V.X.CTRL.TT;
V_D_STEP_shadow <= V.D.STEP;
V_X_CTRL_WICC_shadow <= V.X.CTRL.WICC;
VIR_ADDR31DOWNTO2_shadow <= VIR.ADDR( 31 DOWNTO 2 );
V_M_CTRL_RD7DOWNTO0_shadow <= V.M.CTRL.RD ( 7 DOWNTO 0 );
V_X_RESULT_shadow <= V.X.RESULT;
V_D_CNT_shadow <= V.D.CNT;
XC_VECTT_shadow <= XC_VECTT;
EX_ADD_RES32DOWNTO3_shadow <= EX_ADD_RES ( 32 DOWNTO 3 );
V_W_S_EF_shadow <= V.W.S.EF;
V_A_CTRL_PC31DOWNTO2_shadow <= V.A.CTRL.PC( 31 DOWNTO 2 );
V_X_DATA04DOWNTO0_shadow <= V.X.DATA ( 0 )( 4 DOWNTO 0 );
V_X_DCI_SIGNED_shadow <= V.X.DCI.SIGNED;
V_M_NALIGN_shadow <= V.M.NALIGN;
XC_WREG_shadow <= XC_WREG;
V_A_RFA2_shadow <= V.A.RFA2;
V_E_CTRL_PC31DOWNTO12_shadow <= V.E.CTRL.PC( 31 DOWNTO 12 );
EX_ADD_RES32DOWNTO332DOWNTO13_shadow <= EX_ADD_RES ( 32 DOWNTO 3 )( 32 DOWNTO 13 );
EX_OP231_shadow <= EX_OP2( 31 );
XC_TRAP_ADDRESS31DOWNTO4_shadow <= XC_TRAP_ADDRESS( 31 DOWNTO 4 );
V_X_ICC_shadow <= V.X.ICC;
V_A_SU_shadow <= V.A.SU;
V_E_OP2_shadow <= V.E.OP2;
EX_FORCE_A2_shadow <= EX_FORCE_A2;
V_E_CTRL_PC31DOWNTO2_shadow <= V.E.CTRL.PC( 31 DOWNTO 2 );
V_E_CTRL_PC31DOWNTO4_shadow <= V.E.CTRL.PC( 31 DOWNTO 4 );
V_E_OP131_shadow <= V.E.OP1( 31 );
V_X_DCI_shadow <= V.X.DCI;
V_E_CTRL_WICC_shadow <= V.E.CTRL.WICC;
EX_OP13_shadow <= EX_OP1( 3 );
V_F_PC31DOWNTO12_shadow <= V.F.PC( 31 DOWNTO 12 );
V_E_CTRL_INST_shadow <= V.E.CTRL.INST;
V_E_CTRL_LD_shadow <= V.E.CTRL.LD;
V_M_SU_shadow <= V.M.SU;
V_E_SARI_shadow <= V.E.SARI;
V_E_ET_shadow <= V.E.ET;
V_M_CTRL_PV_shadow <= V.M.CTRL.PV;
VDSU_CRDY2_shadow <= VDSU.CRDY ( 2 );
MUL_OP2_shadow <= MUL_OP2;
XC_EXCEPTION_shadow <= XC_EXCEPTION;
V_E_OP1_shadow <= V.E.OP1;
VP_ERROR_shadow <= VP.ERROR;
V_M_DCI_SIGNED_shadow <= V.M.DCI.SIGNED;
V_D_PC31DOWNTO12_shadow <= V.D.PC( 31 DOWNTO 12 );
MUL_OP231_shadow <= MUL_OP2 ( 31 );
XC_TRAP_ADDRESS31DOWNTO2_shadow <= XC_TRAP_ADDRESS( 31 DOWNTO 2 );
V_M_CTRL_PC3DOWNTO2_shadow <= V.M.CTRL.PC( 3 DOWNTO 2 );
V_M_DCI_shadow <= V.M.DCI;
EX_OP23_shadow <= EX_OP2( 3 );
V_X_CTRL_RD6DOWNTO0_shadow <= V.X.CTRL.RD( 6 DOWNTO 0 );
V_X_CTRL_TRAP_shadow <= V.X.CTRL.TRAP;
V_A_DIVSTART_shadow <= V.A.DIVSTART;
V_X_RESULT6DOWNTO03DOWNTO0_shadow <= V.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 );
VDSU_TT_shadow <= VDSU.TT;
EX_ADD_RES32DOWNTO332DOWNTO5_shadow <= EX_ADD_RES ( 32 DOWNTO 3 )( 32 DOWNTO 5 );
V_X_CTRL_CNT_shadow <= V.X.CTRL.CNT;
V_E_YMSB_shadow <= V.E.YMSB;
EX_ADD_RES32DOWNTO330DOWNTO11_shadow <= EX_ADD_RES ( 32 DOWNTO 3 )( 30 DOWNTO 11 );
V_A_RFE2_shadow <= V.A.RFE2;
V_E_OP13_shadow <= V.E.OP1( 3 );
V_A_CWP_shadow <= V.A.CWP;
ME_SIZE_shadow <= ME_SIZE;
V_X_MAC_shadow <= V.X.MAC;
V_M_CTRL_INST_shadow <= V.M.CTRL.INST;
VIR_ADDR31DOWNTO4_shadow <= VIR.ADDR( 31 DOWNTO 4 );
V_A_CTRL_INST20_shadow <= V.A.CTRL.INST( 20 );
DE_REN2_shadow <= DE_REN2;
V_E_CTRL_PV_shadow <= V.E.CTRL.PV;
V_E_MAC_shadow <= V.E.MAC;
V_X_CTRL_TT3DOWNTO0_shadow <= V.X.CTRL.TT( 3 DOWNTO 0 );
EX_ADD_RES3_shadow <= EX_ADD_RES ( 3 );
V_X_CTRL_INST_shadow <= V.X.CTRL.INST;
V_M_CTRL_PC31DOWNTO2_shadow <= V.M.CTRL.PC( 31 DOWNTO 2 );
V_W_S_ET_shadow <= V.W.S.ET;
V_M_CTRL_CNT_shadow <= V.M.CTRL.CNT;
V_M_CTRL_ANNUL_shadow <= V.M.CTRL.ANNUL;
DE_INST19_shadow <= DE_INST( 19 );
XC_HALT_shadow <= XC_HALT;
V_E_OP231_shadow <= V.E.OP2( 31 );
V_A_CTRL_PC3DOWNTO2_shadow <= V.A.CTRL.PC( 3 DOWNTO 2 );
VIR_ADDR31DOWNTO12_shadow <= VIR.ADDR( 31 DOWNTO 12 );
V_M_CTRL_WICC_shadow <= V.M.CTRL.WICC;
V_M_CTRL_WREG_shadow <= V.M.CTRL.WREG;
V_W_S_S_shadow <= V.W.S.S;
V_F_PC31DOWNTO2_shadow <= V.F.PC( 31 DOWNTO 2 );
V_E_CWP_shadow <= V.E.CWP;
V_A_STEP_shadow <= V.A.STEP;
V_A_CTRL_TT3DOWNTO0_shadow <= V.A.CTRL.TT( 3 DOWNTO 0 );
V_A_CTRL_TRAP_shadow <= V.A.CTRL.TRAP;
NPC31DOWNTO2_shadow <= NPC ( 31 DOWNTO 2 );
V_M_CTRL_TRAP_shadow <= V.M.CTRL.TRAP;
V_D_PC31DOWNTO4_shadow <= V.D.PC( 31 DOWNTO 4 );
V_X_INTACK_shadow <= V.X.INTACK;
SIDLE_shadow <= SIDLE;
V_A_CTRL_RETT_shadow <= V.A.CTRL.RETT;
V_X_DATA03_shadow <= V.X.DATA ( 0 )( 3 );
V_A_CTRL_INST19_shadow <= V.A.CTRL.INST( 19 );
V_W_S_SVT_shadow <= V.W.S.SVT;
V_A_CTRL_PC31DOWNTO4_shadow <= V.A.CTRL.PC( 31 DOWNTO 4 );
V_X_LADDR_shadow <= V.X.LADDR;
V_W_S_DWT_shadow <= V.W.S.DWT;
EX_JUMP_ADDRESS31DOWNTO2_shadow <= EX_JUMP_ADDRESS( 31 DOWNTO 2 );
V_W_S_TBA_shadow <= V.W.S.TBA;
XC_WADDR6DOWNTO0_shadow <= XC_WADDR ( 6 DOWNTO 0 );
V_M_MUL_shadow <= V.M.MUL;
V_E_SU_shadow <= V.E.SU;
V_M_Y31_shadow <= V.M.Y ( 31 );
V_E_OP23_shadow <= V.E.OP2( 3 );
V_M_CTRL_PC31DOWNTO4_shadow <= V.M.CTRL.PC( 31 DOWNTO 4 );
DE_RADDR17DOWNTO0_shadow <= DE_RADDR1 ( 7 DOWNTO 0 );
V_X_CTRL_PC31DOWNTO2_shadow <= V.X.CTRL.PC( 31 DOWNTO 2 );
V_E_CTRL_TRAP_shadow <= V.E.CTRL.TRAP;
V_X_DEBUG_shadow <= V.X.DEBUG;
V_M_DCI_LOCK_shadow <= V.M.DCI.LOCK;
V_X_CTRL_PC3DOWNTO2_shadow <= V.X.CTRL.PC( 3 DOWNTO 2 );
V_X_CTRL_WREG_shadow <= V.X.CTRL.WREG;
V_E_CTRL_INST24_shadow <= V.E.CTRL.INST( 24 );
V_D_MEXC_shadow <= V.D.MEXC;
V_W_RESULT_shadow <= V.W.RESULT;
VFPI_DBG_ENABLE_shadow <= VFPI.DBG.ENABLE;
EX_OP131_shadow <= EX_OP1 ( 31 );
V_D_INST1_shadow <= V.D.INST ( 1 );
V_W_EXCEPT_shadow <= V.W.EXCEPT;
V_E_CTRL_TT3DOWNTO0_shadow <= V.E.CTRL.TT( 3 DOWNTO 0 );
ME_LADDR_shadow <= ME_LADDR;
V_X_CTRL_PC31DOWNTO4_shadow <= V.X.CTRL.PC( 31 DOWNTO 4 );
V_E_CTRL_RETT_shadow <= V.E.CTRL.RETT;
XC_WADDR7DOWNTO0_shadow <= XC_WADDR ( 7 DOWNTO 0 );
V_X_CTRL_PV_shadow <= V.X.CTRL.PV;
V_E_CTRL_RD6DOWNTO0_shadow <= V.E.CTRL.RD( 6 DOWNTO 0 );
V_M_MAC_shadow <= V.M.MAC;
V_D_SET_shadow <= V.D.SET;
VIR_ADDR3DOWNTO2_shadow <= VIR.ADDR( 3 DOWNTO 2 );
V_D_CWP_shadow <= V.D.CWP;
DE_INST20_shadow <= DE_INST( 20 );
V_D_ANNUL_shadow <= V.D.ANNUL;
EX_OP2_shadow <= EX_OP2;
EX_SARI_shadow <= EX_SARI;
V_D_PC31DOWNTO2_shadow <= V.D.PC( 31 DOWNTO 2 );
V_X_DCI_SIZE_shadow <= V.X.DCI.SIZE;
V_M_Y_shadow <= V.M.Y;
V_X_CTRL_PC_shadow <= V.X.CTRL.PC;
V_X_SET_shadow <= V.X.SET;
V_A_CTRL_PC_shadow <= V.A.CTRL.PC;
V_A_JMPL_shadow <= V.A.JMPL;
V_E_CTRL_PC_shadow <= V.E.CTRL.PC;
V_E_CTRL_INST20_shadow <= V.E.CTRL.INST( 20 );
V_E_CTRL_WREG_shadow <= V.E.CTRL.WREG;
V_A_CTRL_WREG_shadow <= V.A.CTRL.WREG;
V_A_CTRL_shadow <= V.A.CTRL;
V_A_CTRL_RD6DOWNTO0_shadow <= V.A.CTRL.RD( 6 DOWNTO 0 );
V_X_DATA0_shadow <= V.X.DATA ( 0 );
V_E_CTRL_INST19_shadow <= V.E.CTRL.INST( 19 );
ME_SIGNED_shadow <= ME_SIGNED;
V_W_WREG_shadow <= V.W.WREG;
V_D_PC_shadow <= V.D.PC;
VFPI_D_ANNUL_shadow <= VFPI.D.ANNUL;
DE_RADDR27DOWNTO0_shadow <= DE_RADDR2 ( 7 DOWNTO 0 );
V_E_CTRL_CNT_shadow <= V.E.CTRL.CNT;
V_F_PC_shadow <= V.F.PC;
V_X_DATA031_shadow <= V.X.DATA ( 0 )( 31 );
V_M_CTRL_PC31DOWNTO12_shadow <= V.M.CTRL.PC( 31 DOWNTO 12 );
V_X_CTRL_RD7DOWNTO0_shadow <= V.X.CTRL.RD ( 7 DOWNTO 0 );
V_M_CTRL_TT_shadow <= V.M.CTRL.TT;
V_X_CTRL_shadow <= V.X.CTRL;
V_A_CTRL_INST24_shadow <= V.A.CTRL.INST( 24 );
XC_TRAP_ADDRESS3DOWNTO2_shadow <= XC_TRAP_ADDRESS( 3 DOWNTO 2 );
V_X_NERROR_shadow <= V.X.NERROR;
V_F_PC31DOWNTO4_shadow <= V.F.PC( 31 DOWNTO 4 );
V_W_S_TT3DOWNTO0_shadow <= V.W.S.TT( 3 DOWNTO 0 );
EX_JUMP_ADDRESS31DOWNTO4_shadow <= EX_JUMP_ADDRESS( 31 DOWNTO 4 );
EX_ADD_RES32DOWNTO332DOWNTO3_shadow <= EX_ADD_RES ( 32 DOWNTO 3 )( 32 DOWNTO 3 );
V_F_BRANCH_shadow <= V.F.BRANCH;
V_A_CTRL_WICC_shadow <= V.A.CTRL.WICC;
V_A_CTRL_LD_shadow <= V.A.CTRL.LD;
V_A_CTRL_TT_shadow <= V.A.CTRL.TT;
V_M_CTRL_LD_shadow <= V.M.CTRL.LD;
V_E_SHCNT_shadow <= V.E.SHCNT;
XC_TRAP_ADDRESS31DOWNTO12_shadow <= XC_TRAP_ADDRESS( 31 DOWNTO 12 );
V_A_CTRL_INST_shadow <= V.A.CTRL.INST;
V_A_CTRL_RD7DOWNTO0_shadow <= V.A.CTRL.RD ( 7 DOWNTO 0 );
VIR_PWD_shadow <= VIR.PWD;
XC_RESULT_shadow <= XC_RESULT;
V_A_RFA1_shadow <= V.A.RFA1;
V_E_JMPL_shadow <= V.E.JMPL;
V_E_CTRL_RD7DOWNTO0_shadow <= V.E.CTRL.RD ( 7 DOWNTO 0 );
ME_ICC_shadow <= ME_ICC;
DE_INST24_shadow <= DE_INST( 24 );
XC_TRAP_shadow <= XC_TRAP;
VDSU_TBUFCNT_shadow <= VDSU.TBUFCNT;
XC_TRAP_ADDRESS_shadow <= XC_TRAP_ADDRESS;
  end process;

dfp_delay : process(clk) begin
	if(clk'event and clk = '1')then
		RPIN_ERROR_intermed_1 <= RPIN.ERROR;
		VP_ERROR_shadow_intermed_1 <= VP_ERROR_shadow;
		V_W_S_S_shadow_intermed_1 <= V_W_S_S_shadow;
		RIN_W_S_S_intermed_1 <= RIN.W.S.S;
		V_W_S_S_shadow_intermed_1 <= V_W_S_S_shadow;
		V_W_S_S_shadow_intermed_2 <= V_W_S_S_shadow_intermed_1;
		V_W_S_PS_shadow_intermed_1 <= V_W_S_PS_shadow;
		RIN_W_S_PS_intermed_1 <= RIN.W.S.PS;
		R_W_S_S_intermed_1 <= R.W.S.S;
		RIN_W_S_S_intermed_1 <= RIN.W.S.S;
		RIN_W_S_S_intermed_2 <= RIN_W_S_S_intermed_1;
		R_X_RESULT6DOWNTO0_intermed_1 <= R.X.RESULT( 6 DOWNTO 0 );
		R_X_RESULT6DOWNTO0_intermed_2 <= R_X_RESULT6DOWNTO0_intermed_1;
		V_X_RESULT6DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO0_shadow;
		V_X_RESULT6DOWNTO0_shadow_intermed_2 <= V_X_RESULT6DOWNTO0_shadow_intermed_1;
		V_X_RESULT6DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO0_shadow;
		RIN_X_RESULT6DOWNTO0_intermed_1 <= RIN.X.RESULT ( 6 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO0_intermed_1 <= RIN.X.RESULT( 6 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO0_intermed_2 <= RIN_X_RESULT6DOWNTO0_intermed_1;
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		V_X_DATA0_shadow_intermed_2 <= V_X_DATA0_shadow_intermed_1;
		R_X_DATA0_intermed_1 <= R.X.DATA( 0 );
		R_X_DATA0_intermed_2 <= R_X_DATA0_intermed_1;
		DCO_DATA0_intermed_1 <= DCO.DATA ( 0 );
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA ( 0 );
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA( 0 );
		RIN_X_DATA0_intermed_2 <= RIN_X_DATA0_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 2 );
		R_M_CTRL_PC31DOWNTO2_intermed_2 <= R_M_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_3 <= RIN_M_CTRL_PC31DOWNTO2_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		RIN_A_CTRL_PC31DOWNTO2_intermed_5 <= RIN_A_CTRL_PC31DOWNTO2_intermed_4;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_4 <= R_A_CTRL_PC31DOWNTO2_intermed_3;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC ( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		R_X_CTRL_PC31DOWNTO2_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 2 );
		R_X_CTRL_PC31DOWNTO2_intermed_2 <= R_X_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC ( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_5 <= V_D_PC31DOWNTO2_shadow_intermed_4;
		V_D_PC31DOWNTO2_shadow_intermed_6 <= V_D_PC31DOWNTO2_shadow_intermed_5;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_5 <= RIN_D_PC31DOWNTO2_intermed_4;
		RIN_D_PC31DOWNTO2_intermed_6 <= RIN_D_PC31DOWNTO2_intermed_5;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC ( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC ( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC ( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_2 <= RIN_X_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC ( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_3 <= R_E_CTRL_PC31DOWNTO2_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		R_D_PC31DOWNTO2_intermed_4 <= R_D_PC31DOWNTO2_intermed_3;
		R_D_PC31DOWNTO2_intermed_5 <= R_D_PC31DOWNTO2_intermed_4;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC ( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_4 <= RIN_E_CTRL_PC31DOWNTO2_intermed_3;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO2_shadow;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_X_ANNUL_ALL_shadow_intermed_1 <= V_X_ANNUL_ALL_shadow;
		V_X_ANNUL_ALL_shadow_intermed_2 <= V_X_ANNUL_ALL_shadow_intermed_1;
		V_X_ANNUL_ALL_shadow_intermed_3 <= V_X_ANNUL_ALL_shadow_intermed_2;
		V_X_ANNUL_ALL_shadow_intermed_4 <= V_X_ANNUL_ALL_shadow_intermed_3;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_A_CTRL_ANNUL_intermed_2 <= RIN_A_CTRL_ANNUL_intermed_1;
		RIN_A_CTRL_ANNUL_intermed_3 <= RIN_A_CTRL_ANNUL_intermed_2;
		RIN_A_CTRL_ANNUL_intermed_4 <= RIN_A_CTRL_ANNUL_intermed_3;
		RIN_A_CTRL_ANNUL_intermed_5 <= RIN_A_CTRL_ANNUL_intermed_4;
		R_M_CTRL_WREG_intermed_1 <= R.M.CTRL.WREG;
		R_A_CTRL_ANNUL_intermed_1 <= R.A.CTRL.ANNUL;
		R_A_CTRL_ANNUL_intermed_2 <= R_A_CTRL_ANNUL_intermed_1;
		R_A_CTRL_ANNUL_intermed_3 <= R_A_CTRL_ANNUL_intermed_2;
		R_A_CTRL_ANNUL_intermed_4 <= R_A_CTRL_ANNUL_intermed_3;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_X_ANNUL_ALL_intermed_2 <= RIN_X_ANNUL_ALL_intermed_1;
		RIN_X_ANNUL_ALL_intermed_3 <= RIN_X_ANNUL_ALL_intermed_2;
		RIN_X_ANNUL_ALL_intermed_4 <= RIN_X_ANNUL_ALL_intermed_3;
		RIN_X_ANNUL_ALL_intermed_5 <= RIN_X_ANNUL_ALL_intermed_4;
		V_M_CTRL_WREG_shadow_intermed_1 <= V_M_CTRL_WREG_shadow;
		V_M_CTRL_WREG_shadow_intermed_2 <= V_M_CTRL_WREG_shadow_intermed_1;
		R_X_ANNUL_ALL_intermed_1 <= R.X.ANNUL_ALL;
		R_X_ANNUL_ALL_intermed_2 <= R_X_ANNUL_ALL_intermed_1;
		R_X_ANNUL_ALL_intermed_3 <= R_X_ANNUL_ALL_intermed_2;
		R_X_ANNUL_ALL_intermed_4 <= R_X_ANNUL_ALL_intermed_3;
		V_X_CTRL_WREG_shadow_intermed_1 <= V_X_CTRL_WREG_shadow;
		R_E_CTRL_WREG_intermed_1 <= R.E.CTRL.WREG;
		R_E_CTRL_WREG_intermed_2 <= R_E_CTRL_WREG_intermed_1;
		RIN_X_CTRL_WREG_intermed_1 <= RIN.X.CTRL.WREG;
		V_A_CTRL_ANNUL_shadow_intermed_1 <= V_A_CTRL_ANNUL_shadow;
		V_A_CTRL_ANNUL_shadow_intermed_2 <= V_A_CTRL_ANNUL_shadow_intermed_1;
		V_A_CTRL_ANNUL_shadow_intermed_3 <= V_A_CTRL_ANNUL_shadow_intermed_2;
		V_A_CTRL_ANNUL_shadow_intermed_4 <= V_A_CTRL_ANNUL_shadow_intermed_3;
		RIN_E_CTRL_WREG_intermed_1 <= RIN.E.CTRL.WREG;
		RIN_E_CTRL_WREG_intermed_2 <= RIN_E_CTRL_WREG_intermed_1;
		RIN_E_CTRL_WREG_intermed_3 <= RIN_E_CTRL_WREG_intermed_2;
		RIN_M_CTRL_WREG_intermed_1 <= RIN.M.CTRL.WREG;
		RIN_M_CTRL_WREG_intermed_2 <= RIN_M_CTRL_WREG_intermed_1;
		V_E_CTRL_WREG_shadow_intermed_1 <= V_E_CTRL_WREG_shadow;
		V_E_CTRL_WREG_shadow_intermed_2 <= V_E_CTRL_WREG_shadow_intermed_1;
		V_E_CTRL_WREG_shadow_intermed_3 <= V_E_CTRL_WREG_shadow_intermed_2;
		RIN_A_CTRL_WREG_intermed_1 <= RIN.A.CTRL.WREG;
		RIN_A_CTRL_WREG_intermed_2 <= RIN_A_CTRL_WREG_intermed_1;
		RIN_A_CTRL_WREG_intermed_3 <= RIN_A_CTRL_WREG_intermed_2;
		RIN_A_CTRL_WREG_intermed_4 <= RIN_A_CTRL_WREG_intermed_3;
		V_A_CTRL_WREG_shadow_intermed_1 <= V_A_CTRL_WREG_shadow;
		V_A_CTRL_WREG_shadow_intermed_2 <= V_A_CTRL_WREG_shadow_intermed_1;
		V_A_CTRL_WREG_shadow_intermed_3 <= V_A_CTRL_WREG_shadow_intermed_2;
		V_A_CTRL_WREG_shadow_intermed_4 <= V_A_CTRL_WREG_shadow_intermed_3;
		R_A_CTRL_WREG_intermed_1 <= R.A.CTRL.WREG;
		R_A_CTRL_WREG_intermed_2 <= R_A_CTRL_WREG_intermed_1;
		R_A_CTRL_WREG_intermed_3 <= R_A_CTRL_WREG_intermed_2;
		RIN_X_INTACK_intermed_1 <= RIN.X.INTACK;
		V_X_INTACK_shadow_intermed_1 <= V_X_INTACK_shadow;
		V_X_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_X_CTRL_TT3DOWNTO0_shadow;
		V_X_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_X_CTRL_TT3DOWNTO0_shadow_intermed_1;
		V_X_CTRL_TT3DOWNTO0_shadow_intermed_3 <= V_X_CTRL_TT3DOWNTO0_shadow_intermed_2;
		R_M_CTRL_TT3DOWNTO0_intermed_1 <= R.M.CTRL.TT( 3 DOWNTO 0 );
		R_M_CTRL_TT3DOWNTO0_intermed_2 <= R_M_CTRL_TT3DOWNTO0_intermed_1;
		R_M_CTRL_TT3DOWNTO0_intermed_3 <= R_M_CTRL_TT3DOWNTO0_intermed_2;
		V_M_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_M_CTRL_TT3DOWNTO0_shadow;
		V_M_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_M_CTRL_TT3DOWNTO0_shadow_intermed_1;
		V_M_CTRL_TT3DOWNTO0_shadow_intermed_3 <= V_M_CTRL_TT3DOWNTO0_shadow_intermed_2;
		V_M_CTRL_TT3DOWNTO0_shadow_intermed_4 <= V_M_CTRL_TT3DOWNTO0_shadow_intermed_3;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_3 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_4 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_3;
		R_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= R.X.RESULT( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		R_X_RESULT6DOWNTO03DOWNTO0_intermed_2 <= R_X_RESULT6DOWNTO03DOWNTO0_intermed_1;
		R_X_RESULT6DOWNTO03DOWNTO0_intermed_3 <= R_X_RESULT6DOWNTO03DOWNTO0_intermed_2;
		R_A_CTRL_TT3DOWNTO0_intermed_1 <= R.A.CTRL.TT( 3 DOWNTO 0 );
		R_A_CTRL_TT3DOWNTO0_intermed_2 <= R_A_CTRL_TT3DOWNTO0_intermed_1;
		R_A_CTRL_TT3DOWNTO0_intermed_3 <= R_A_CTRL_TT3DOWNTO0_intermed_2;
		R_A_CTRL_TT3DOWNTO0_intermed_4 <= R_A_CTRL_TT3DOWNTO0_intermed_3;
		R_A_CTRL_TT3DOWNTO0_intermed_5 <= R_A_CTRL_TT3DOWNTO0_intermed_4;
		RIN_A_CTRL_TT3DOWNTO0_intermed_1 <= RIN.A.CTRL.TT( 3 DOWNTO 0 );
		RIN_A_CTRL_TT3DOWNTO0_intermed_2 <= RIN_A_CTRL_TT3DOWNTO0_intermed_1;
		RIN_A_CTRL_TT3DOWNTO0_intermed_3 <= RIN_A_CTRL_TT3DOWNTO0_intermed_2;
		RIN_A_CTRL_TT3DOWNTO0_intermed_4 <= RIN_A_CTRL_TT3DOWNTO0_intermed_3;
		RIN_A_CTRL_TT3DOWNTO0_intermed_5 <= RIN_A_CTRL_TT3DOWNTO0_intermed_4;
		RIN_A_CTRL_TT3DOWNTO0_intermed_6 <= RIN_A_CTRL_TT3DOWNTO0_intermed_5;
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= RIN.X.RESULT( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2 <= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1;
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_3 <= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2;
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_4 <= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_3;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_A_CTRL_TT3DOWNTO0_shadow;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_1;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_3 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_2;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_4 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_3;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_5 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_4;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_6 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_5;
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= RIN.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2 <= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1;
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_3 <= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2;
		R_W_S_TT3DOWNTO0_intermed_1 <= R.W.S.TT( 3 DOWNTO 0 );
		R_W_S_TT3DOWNTO0_intermed_2 <= R_W_S_TT3DOWNTO0_intermed_1;
		R_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= R.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		R_X_RESULT6DOWNTO03DOWNTO0_intermed_2 <= R_X_RESULT6DOWNTO03DOWNTO0_intermed_1;
		R_E_CTRL_TT3DOWNTO0_intermed_1 <= R.E.CTRL.TT( 3 DOWNTO 0 );
		R_E_CTRL_TT3DOWNTO0_intermed_2 <= R_E_CTRL_TT3DOWNTO0_intermed_1;
		R_E_CTRL_TT3DOWNTO0_intermed_3 <= R_E_CTRL_TT3DOWNTO0_intermed_2;
		R_E_CTRL_TT3DOWNTO0_intermed_4 <= R_E_CTRL_TT3DOWNTO0_intermed_3;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_3 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2;
		RIN_W_S_TT3DOWNTO0_intermed_1 <= RIN.W.S.TT( 3 DOWNTO 0 );
		RIN_W_S_TT3DOWNTO0_intermed_2 <= RIN_W_S_TT3DOWNTO0_intermed_1;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_E_CTRL_TT3DOWNTO0_shadow;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_E_CTRL_TT3DOWNTO0_shadow_intermed_1;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_3 <= V_E_CTRL_TT3DOWNTO0_shadow_intermed_2;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_4 <= V_E_CTRL_TT3DOWNTO0_shadow_intermed_3;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_5 <= V_E_CTRL_TT3DOWNTO0_shadow_intermed_4;
		RIN_W_S_TT3DOWNTO0_intermed_1 <= RIN.W.S.TT ( 3 DOWNTO 0 );
		RIN_M_CTRL_TT3DOWNTO0_intermed_1 <= RIN.M.CTRL.TT( 3 DOWNTO 0 );
		RIN_M_CTRL_TT3DOWNTO0_intermed_2 <= RIN_M_CTRL_TT3DOWNTO0_intermed_1;
		RIN_M_CTRL_TT3DOWNTO0_intermed_3 <= RIN_M_CTRL_TT3DOWNTO0_intermed_2;
		RIN_M_CTRL_TT3DOWNTO0_intermed_4 <= RIN_M_CTRL_TT3DOWNTO0_intermed_3;
		RIN_X_CTRL_TT3DOWNTO0_intermed_1 <= RIN.X.CTRL.TT( 3 DOWNTO 0 );
		RIN_X_CTRL_TT3DOWNTO0_intermed_2 <= RIN_X_CTRL_TT3DOWNTO0_intermed_1;
		RIN_X_CTRL_TT3DOWNTO0_intermed_3 <= RIN_X_CTRL_TT3DOWNTO0_intermed_2;
		V_W_S_TT3DOWNTO0_shadow_intermed_1 <= V_W_S_TT3DOWNTO0_shadow;
		V_W_S_TT3DOWNTO0_shadow_intermed_2 <= V_W_S_TT3DOWNTO0_shadow_intermed_1;
		R_X_CTRL_TT3DOWNTO0_intermed_1 <= R.X.CTRL.TT( 3 DOWNTO 0 );
		R_X_CTRL_TT3DOWNTO0_intermed_2 <= R_X_CTRL_TT3DOWNTO0_intermed_1;
		RIN_E_CTRL_TT3DOWNTO0_intermed_1 <= RIN.E.CTRL.TT( 3 DOWNTO 0 );
		RIN_E_CTRL_TT3DOWNTO0_intermed_2 <= RIN_E_CTRL_TT3DOWNTO0_intermed_1;
		RIN_E_CTRL_TT3DOWNTO0_intermed_3 <= RIN_E_CTRL_TT3DOWNTO0_intermed_2;
		RIN_E_CTRL_TT3DOWNTO0_intermed_4 <= RIN_E_CTRL_TT3DOWNTO0_intermed_3;
		RIN_E_CTRL_TT3DOWNTO0_intermed_5 <= RIN_E_CTRL_TT3DOWNTO0_intermed_4;
		V_W_S_TT3DOWNTO0_shadow_intermed_1 <= V_W_S_TT3DOWNTO0_shadow;
		XC_VECTT3DOWNTO0_shadow_intermed_1 <= XC_VECTT3DOWNTO0_shadow;
		XC_VECTT3DOWNTO0_shadow_intermed_2 <= XC_VECTT3DOWNTO0_shadow_intermed_1;
		RIN_X_INTACK_intermed_1 <= RIN.X.INTACK;
		V_X_INTACK_shadow_intermed_1 <= V_X_INTACK_shadow;
		V_M_RESULT1DOWNTO0_shadow_intermed_1 <= V_M_RESULT1DOWNTO0_shadow;
		V_M_RESULT1DOWNTO0_shadow_intermed_2 <= V_M_RESULT1DOWNTO0_shadow_intermed_1;
		RIN_M_RESULT1DOWNTO0_intermed_1 <= RIN.M.RESULT ( 1 DOWNTO 0 );
		RIN_M_RESULT1DOWNTO0_intermed_1 <= RIN.M.RESULT( 1 DOWNTO 0 );
		RIN_M_RESULT1DOWNTO0_intermed_2 <= RIN_M_RESULT1DOWNTO0_intermed_1;
		V_M_RESULT1DOWNTO0_shadow_intermed_1 <= V_M_RESULT1DOWNTO0_shadow;
		R_M_RESULT1DOWNTO0_intermed_1 <= R.M.RESULT( 1 DOWNTO 0 );
		R_M_RESULT1DOWNTO0_intermed_2 <= R_M_RESULT1DOWNTO0_intermed_1;
		V_X_ANNUL_ALL_shadow_intermed_1 <= V_X_ANNUL_ALL_shadow;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_A_CTRL_ANNUL_intermed_2 <= RIN_A_CTRL_ANNUL_intermed_1;
		RIN_A_CTRL_ANNUL_intermed_3 <= RIN_A_CTRL_ANNUL_intermed_2;
		RIN_E_CTRL_ANNUL_intermed_1 <= RIN.E.CTRL.ANNUL;
		RIN_E_CTRL_ANNUL_intermed_2 <= RIN_E_CTRL_ANNUL_intermed_1;
		R_A_CTRL_ANNUL_intermed_1 <= R.A.CTRL.ANNUL;
		R_A_CTRL_ANNUL_intermed_2 <= R_A_CTRL_ANNUL_intermed_1;
		V_M_CTRL_ANNUL_shadow_intermed_1 <= V_M_CTRL_ANNUL_shadow;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_X_ANNUL_ALL_intermed_2 <= RIN_X_ANNUL_ALL_intermed_1;
		R_X_ANNUL_ALL_intermed_1 <= R.X.ANNUL_ALL;
		RIN_M_DCI_LOCK_intermed_1 <= RIN.M.DCI.LOCK;
		V_E_CTRL_ANNUL_shadow_intermed_1 <= V_E_CTRL_ANNUL_shadow;
		V_E_CTRL_ANNUL_shadow_intermed_2 <= V_E_CTRL_ANNUL_shadow_intermed_1;
		V_A_CTRL_ANNUL_shadow_intermed_1 <= V_A_CTRL_ANNUL_shadow;
		V_A_CTRL_ANNUL_shadow_intermed_2 <= V_A_CTRL_ANNUL_shadow_intermed_1;
		V_A_CTRL_ANNUL_shadow_intermed_3 <= V_A_CTRL_ANNUL_shadow_intermed_2;
		RIN_M_CTRL_ANNUL_intermed_1 <= RIN.M.CTRL.ANNUL;
		R_E_CTRL_ANNUL_intermed_1 <= R.E.CTRL.ANNUL;
		V_M_DCI_LOCK_shadow_intermed_1 <= V_M_DCI_LOCK_shadow;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA ( 0 )( 31 );
		RIN_X_DATA031_intermed_2 <= RIN_X_DATA031_intermed_1;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_2 <= V_X_DATA031_shadow_intermed_1;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_2 <= V_X_DATA031_shadow_intermed_1;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA( 0 )( 31 );
		RIN_X_DATA031_intermed_2 <= RIN_X_DATA031_intermed_1;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA ( 0 ) ( 31 );
		DCO_DATA031_intermed_1 <= DCO.DATA ( 0 )( 31 );
		DCO_DATA031_intermed_2 <= DCO_DATA031_intermed_1;
		R_X_DATA031_intermed_1 <= R.X.DATA( 0 )( 31 );
		R_X_DATA031_intermed_2 <= R_X_DATA031_intermed_1;
		R_X_DATA031_intermed_1 <= R.X.DATA ( 0 )( 31 );
		R_X_DATA031_intermed_2 <= R_X_DATA031_intermed_1;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		DE_INST19_shadow_intermed_1 <= DE_INST19_shadow;
		DE_INST19_shadow_intermed_2 <= DE_INST19_shadow_intermed_1;
		DE_INST19_shadow_intermed_3 <= DE_INST19_shadow_intermed_2;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_3 <= V_A_CTRL_INST19_shadow_intermed_2;
		V_E_CTRL_INST19_shadow_intermed_1 <= V_E_CTRL_INST19_shadow;
		V_E_CTRL_INST19_shadow_intermed_1 <= V_E_CTRL_INST19_shadow;
		V_E_CTRL_INST19_shadow_intermed_2 <= V_E_CTRL_INST19_shadow_intermed_1;
		R_E_CTRL_INST19_intermed_1 <= R.E.CTRL.INST( 19 );
		R_E_CTRL_INST19_intermed_2 <= R_E_CTRL_INST19_intermed_1;
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST ( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST( 19 );
		R_A_CTRL_INST19_intermed_2 <= R_A_CTRL_INST19_intermed_1;
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST ( 19 );
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		RIN_A_CTRL_INST19_intermed_3 <= RIN_A_CTRL_INST19_intermed_2;
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST ( 19 );
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST( 19 );
		RIN_E_CTRL_INST19_intermed_2 <= RIN_E_CTRL_INST19_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		V_A_CTRL_INST20_shadow_intermed_1 <= V_A_CTRL_INST20_shadow;
		V_A_CTRL_INST20_shadow_intermed_2 <= V_A_CTRL_INST20_shadow_intermed_1;
		RIN_A_CTRL_INST20_intermed_1 <= RIN.A.CTRL.INST ( 20 );
		RIN_A_CTRL_INST20_intermed_2 <= RIN_A_CTRL_INST20_intermed_1;
		RIN_E_CTRL_INST20_intermed_1 <= RIN.E.CTRL.INST ( 20 );
		R_A_CTRL_INST20_intermed_1 <= R.A.CTRL.INST ( 20 );
		R_E_CTRL_INST20_intermed_1 <= R.E.CTRL.INST( 20 );
		R_E_CTRL_INST20_intermed_2 <= R_E_CTRL_INST20_intermed_1;
		RIN_A_CTRL_INST20_intermed_1 <= RIN.A.CTRL.INST( 20 );
		RIN_A_CTRL_INST20_intermed_2 <= RIN_A_CTRL_INST20_intermed_1;
		RIN_A_CTRL_INST20_intermed_3 <= RIN_A_CTRL_INST20_intermed_2;
		V_E_CTRL_INST20_shadow_intermed_1 <= V_E_CTRL_INST20_shadow;
		V_E_CTRL_INST20_shadow_intermed_2 <= V_E_CTRL_INST20_shadow_intermed_1;
		V_E_CTRL_INST20_shadow_intermed_1 <= V_E_CTRL_INST20_shadow;
		DE_INST20_shadow_intermed_1 <= DE_INST20_shadow;
		DE_INST20_shadow_intermed_2 <= DE_INST20_shadow_intermed_1;
		DE_INST20_shadow_intermed_3 <= DE_INST20_shadow_intermed_2;
		V_A_CTRL_INST20_shadow_intermed_1 <= V_A_CTRL_INST20_shadow;
		V_A_CTRL_INST20_shadow_intermed_2 <= V_A_CTRL_INST20_shadow_intermed_1;
		V_A_CTRL_INST20_shadow_intermed_3 <= V_A_CTRL_INST20_shadow_intermed_2;
		RIN_E_CTRL_INST20_intermed_1 <= RIN.E.CTRL.INST( 20 );
		RIN_E_CTRL_INST20_intermed_2 <= RIN_E_CTRL_INST20_intermed_1;
		R_A_CTRL_INST20_intermed_1 <= R.A.CTRL.INST( 20 );
		R_A_CTRL_INST20_intermed_2 <= R_A_CTRL_INST20_intermed_1;
		RIN_X_DATA00_intermed_1 <= RIN.X.DATA ( 0 )( 0 );
		RIN_X_DATA00_intermed_2 <= RIN_X_DATA00_intermed_1;
		V_X_DATA00_shadow_intermed_1 <= V_X_DATA00_shadow;
		DCO_DATA00_intermed_1 <= DCO.DATA ( 0 )( 0 );
		DCO_DATA00_intermed_2 <= DCO_DATA00_intermed_1;
		V_X_DATA00_shadow_intermed_1 <= V_X_DATA00_shadow;
		V_X_DATA00_shadow_intermed_2 <= V_X_DATA00_shadow_intermed_1;
		RIN_X_DATA00_intermed_1 <= RIN.X.DATA ( 0 ) ( 0 );
		V_X_DATA00_shadow_intermed_1 <= V_X_DATA00_shadow;
		V_X_DATA00_shadow_intermed_2 <= V_X_DATA00_shadow_intermed_1;
		R_X_DATA00_intermed_1 <= R.X.DATA ( 0 )( 0 );
		R_X_DATA00_intermed_2 <= R_X_DATA00_intermed_1;
		RIN_X_DATA00_intermed_1 <= RIN.X.DATA( 0 )( 0 );
		RIN_X_DATA00_intermed_2 <= RIN_X_DATA00_intermed_1;
		R_X_DATA00_intermed_1 <= R.X.DATA( 0 )( 0 );
		R_X_DATA00_intermed_2 <= R_X_DATA00_intermed_1;
		RIN_X_DATA04DOWNTO0_intermed_1 <= RIN.X.DATA ( 0 ) ( 4 DOWNTO 0 );
		V_X_DATA04DOWNTO0_shadow_intermed_1 <= V_X_DATA04DOWNTO0_shadow;
		V_X_DATA04DOWNTO0_shadow_intermed_2 <= V_X_DATA04DOWNTO0_shadow_intermed_1;
		R_X_DATA04DOWNTO0_intermed_1 <= R.X.DATA( 0 )( 4 DOWNTO 0 );
		R_X_DATA04DOWNTO0_intermed_2 <= R_X_DATA04DOWNTO0_intermed_1;
		R_X_DATA04DOWNTO0_intermed_1 <= R.X.DATA ( 0 )( 4 DOWNTO 0 );
		R_X_DATA04DOWNTO0_intermed_2 <= R_X_DATA04DOWNTO0_intermed_1;
		V_X_DATA04DOWNTO0_shadow_intermed_1 <= V_X_DATA04DOWNTO0_shadow;
		DCO_DATA04DOWNTO0_intermed_1 <= DCO.DATA ( 0 )( 4 DOWNTO 0 );
		DCO_DATA04DOWNTO0_intermed_2 <= DCO_DATA04DOWNTO0_intermed_1;
		RIN_X_DATA04DOWNTO0_intermed_1 <= RIN.X.DATA ( 0 )( 4 DOWNTO 0 );
		RIN_X_DATA04DOWNTO0_intermed_2 <= RIN_X_DATA04DOWNTO0_intermed_1;
		RIN_X_DATA04DOWNTO0_intermed_1 <= RIN.X.DATA( 0 )( 4 DOWNTO 0 );
		RIN_X_DATA04DOWNTO0_intermed_2 <= RIN_X_DATA04DOWNTO0_intermed_1;
		V_X_DATA04DOWNTO0_shadow_intermed_1 <= V_X_DATA04DOWNTO0_shadow;
		V_X_DATA04DOWNTO0_shadow_intermed_2 <= V_X_DATA04DOWNTO0_shadow_intermed_1;
		RIN_A_RFE1_intermed_1 <= RIN.A.RFE1;
		V_A_RFE1_shadow_intermed_1 <= V_A_RFE1_shadow;
		RIN_A_RFE2_intermed_1 <= RIN.A.RFE2;
		V_A_RFE2_shadow_intermed_1 <= V_A_RFE2_shadow;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 2 );
		R_M_CTRL_PC31DOWNTO2_intermed_2 <= R_M_CTRL_PC31DOWNTO2_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_3 <= R_M_CTRL_PC31DOWNTO2_intermed_2;
		R_M_CTRL_PC31DOWNTO2_intermed_4 <= R_M_CTRL_PC31DOWNTO2_intermed_3;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_3 <= RIN_M_CTRL_PC31DOWNTO2_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_4 <= RIN_M_CTRL_PC31DOWNTO2_intermed_3;
		RIN_M_CTRL_PC31DOWNTO2_intermed_5 <= RIN_M_CTRL_PC31DOWNTO2_intermed_4;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_4;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_6 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_5;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		RIN_A_CTRL_PC31DOWNTO2_intermed_5 <= RIN_A_CTRL_PC31DOWNTO2_intermed_4;
		RIN_A_CTRL_PC31DOWNTO2_intermed_6 <= RIN_A_CTRL_PC31DOWNTO2_intermed_5;
		RIN_A_CTRL_PC31DOWNTO2_intermed_7 <= RIN_A_CTRL_PC31DOWNTO2_intermed_6;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_4 <= R_A_CTRL_PC31DOWNTO2_intermed_3;
		R_A_CTRL_PC31DOWNTO2_intermed_5 <= R_A_CTRL_PC31DOWNTO2_intermed_4;
		R_A_CTRL_PC31DOWNTO2_intermed_6 <= R_A_CTRL_PC31DOWNTO2_intermed_5;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_4;
		R_X_CTRL_PC31DOWNTO2_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 2 );
		R_X_CTRL_PC31DOWNTO2_intermed_2 <= R_X_CTRL_PC31DOWNTO2_intermed_1;
		R_X_CTRL_PC31DOWNTO2_intermed_3 <= R_X_CTRL_PC31DOWNTO2_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_5 <= V_D_PC31DOWNTO2_shadow_intermed_4;
		V_D_PC31DOWNTO2_shadow_intermed_6 <= V_D_PC31DOWNTO2_shadow_intermed_5;
		V_D_PC31DOWNTO2_shadow_intermed_7 <= V_D_PC31DOWNTO2_shadow_intermed_6;
		V_D_PC31DOWNTO2_shadow_intermed_8 <= V_D_PC31DOWNTO2_shadow_intermed_7;
		XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_1 <= XC_TRAP_ADDRESS31DOWNTO2_shadow;
		XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_2 <= XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_5 <= RIN_D_PC31DOWNTO2_intermed_4;
		RIN_D_PC31DOWNTO2_intermed_6 <= RIN_D_PC31DOWNTO2_intermed_5;
		RIN_D_PC31DOWNTO2_intermed_7 <= RIN_D_PC31DOWNTO2_intermed_6;
		RIN_D_PC31DOWNTO2_intermed_8 <= RIN_D_PC31DOWNTO2_intermed_7;
		EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_1 <= EX_ADD_RES32DOWNTO332DOWNTO3_shadow;
		EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_2 <= EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_1;
		V_F_PC31DOWNTO2_shadow_intermed_1 <= V_F_PC31DOWNTO2_shadow;
		V_F_PC31DOWNTO2_shadow_intermed_2 <= V_F_PC31DOWNTO2_shadow_intermed_1;
		V_F_PC31DOWNTO2_shadow_intermed_1 <= V_F_PC31DOWNTO2_shadow;
		RIN_F_PC31DOWNTO2_intermed_1 <= RIN.F.PC( 31 DOWNTO 2 );
		RIN_F_PC31DOWNTO2_intermed_2 <= RIN_F_PC31DOWNTO2_intermed_1;
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_2 <= RIN_X_CTRL_PC31DOWNTO2_intermed_1;
		RIN_X_CTRL_PC31DOWNTO2_intermed_3 <= RIN_X_CTRL_PC31DOWNTO2_intermed_2;
		RIN_X_CTRL_PC31DOWNTO2_intermed_4 <= RIN_X_CTRL_PC31DOWNTO2_intermed_3;
		IRIN_ADDR31DOWNTO2_intermed_1 <= IRIN.ADDR( 31 DOWNTO 2 );
		IRIN_ADDR31DOWNTO2_intermed_2 <= IRIN_ADDR31DOWNTO2_intermed_1;
		IRIN_ADDR31DOWNTO2_intermed_3 <= IRIN_ADDR31DOWNTO2_intermed_2;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_3 <= R_E_CTRL_PC31DOWNTO2_intermed_2;
		R_E_CTRL_PC31DOWNTO2_intermed_4 <= R_E_CTRL_PC31DOWNTO2_intermed_3;
		R_E_CTRL_PC31DOWNTO2_intermed_5 <= R_E_CTRL_PC31DOWNTO2_intermed_4;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_6 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_5;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_7 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_6;
		EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_1 <= EX_JUMP_ADDRESS31DOWNTO2_shadow;
		EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_2 <= EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_1;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		R_D_PC31DOWNTO2_intermed_4 <= R_D_PC31DOWNTO2_intermed_3;
		R_D_PC31DOWNTO2_intermed_5 <= R_D_PC31DOWNTO2_intermed_4;
		R_D_PC31DOWNTO2_intermed_6 <= R_D_PC31DOWNTO2_intermed_5;
		R_D_PC31DOWNTO2_intermed_7 <= R_D_PC31DOWNTO2_intermed_6;
		RIN_F_PC31DOWNTO2_intermed_1 <= RIN.F.PC ( 31 DOWNTO 2 );
		IR_ADDR31DOWNTO2_intermed_1 <= IR.ADDR( 31 DOWNTO 2 );
		IR_ADDR31DOWNTO2_intermed_2 <= IR_ADDR31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_4 <= RIN_E_CTRL_PC31DOWNTO2_intermed_3;
		RIN_E_CTRL_PC31DOWNTO2_intermed_5 <= RIN_E_CTRL_PC31DOWNTO2_intermed_4;
		RIN_E_CTRL_PC31DOWNTO2_intermed_6 <= RIN_E_CTRL_PC31DOWNTO2_intermed_5;
		R_F_PC31DOWNTO2_intermed_1 <= R.F.PC( 31 DOWNTO 2 );
		R_F_PC31DOWNTO2_intermed_2 <= R_F_PC31DOWNTO2_intermed_1;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO2_shadow;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_3;
		VIR_ADDR31DOWNTO2_shadow_intermed_1 <= VIR_ADDR31DOWNTO2_shadow;
		VIR_ADDR31DOWNTO2_shadow_intermed_2 <= VIR_ADDR31DOWNTO2_shadow_intermed_1;
		VIR_ADDR31DOWNTO2_shadow_intermed_3 <= VIR_ADDR31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC ( 31 DOWNTO 2 );
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC ( 31 DOWNTO 2 );
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 2 );
		R_M_CTRL_PC31DOWNTO2_intermed_2 <= R_M_CTRL_PC31DOWNTO2_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_3 <= R_M_CTRL_PC31DOWNTO2_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_3 <= RIN_M_CTRL_PC31DOWNTO2_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_4 <= RIN_M_CTRL_PC31DOWNTO2_intermed_3;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_4;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		RIN_A_CTRL_PC31DOWNTO2_intermed_5 <= RIN_A_CTRL_PC31DOWNTO2_intermed_4;
		RIN_A_CTRL_PC31DOWNTO2_intermed_6 <= RIN_A_CTRL_PC31DOWNTO2_intermed_5;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_4 <= R_A_CTRL_PC31DOWNTO2_intermed_3;
		R_A_CTRL_PC31DOWNTO2_intermed_5 <= R_A_CTRL_PC31DOWNTO2_intermed_4;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_3;
		R_X_CTRL_PC31DOWNTO2_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 2 );
		R_X_CTRL_PC31DOWNTO2_intermed_2 <= R_X_CTRL_PC31DOWNTO2_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_5 <= V_D_PC31DOWNTO2_shadow_intermed_4;
		V_D_PC31DOWNTO2_shadow_intermed_6 <= V_D_PC31DOWNTO2_shadow_intermed_5;
		V_D_PC31DOWNTO2_shadow_intermed_7 <= V_D_PC31DOWNTO2_shadow_intermed_6;
		XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_1 <= XC_TRAP_ADDRESS31DOWNTO2_shadow;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_5 <= RIN_D_PC31DOWNTO2_intermed_4;
		RIN_D_PC31DOWNTO2_intermed_6 <= RIN_D_PC31DOWNTO2_intermed_5;
		RIN_D_PC31DOWNTO2_intermed_7 <= RIN_D_PC31DOWNTO2_intermed_6;
		EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_1 <= EX_ADD_RES32DOWNTO332DOWNTO3_shadow;
		EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_2 <= EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_1;
		V_F_PC31DOWNTO2_shadow_intermed_1 <= V_F_PC31DOWNTO2_shadow;
		V_F_PC31DOWNTO2_shadow_intermed_2 <= V_F_PC31DOWNTO2_shadow_intermed_1;
		V_F_PC31DOWNTO2_shadow_intermed_1 <= V_F_PC31DOWNTO2_shadow;
		RIN_F_PC31DOWNTO2_intermed_1 <= RIN.F.PC( 31 DOWNTO 2 );
		RIN_F_PC31DOWNTO2_intermed_2 <= RIN_F_PC31DOWNTO2_intermed_1;
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_2 <= RIN_X_CTRL_PC31DOWNTO2_intermed_1;
		RIN_X_CTRL_PC31DOWNTO2_intermed_3 <= RIN_X_CTRL_PC31DOWNTO2_intermed_2;
		IRIN_ADDR31DOWNTO2_intermed_1 <= IRIN.ADDR( 31 DOWNTO 2 );
		IRIN_ADDR31DOWNTO2_intermed_2 <= IRIN_ADDR31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_3 <= R_E_CTRL_PC31DOWNTO2_intermed_2;
		R_E_CTRL_PC31DOWNTO2_intermed_4 <= R_E_CTRL_PC31DOWNTO2_intermed_3;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_6 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_5;
		EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_1 <= EX_JUMP_ADDRESS31DOWNTO2_shadow;
		EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_2 <= EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_1;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		R_D_PC31DOWNTO2_intermed_4 <= R_D_PC31DOWNTO2_intermed_3;
		R_D_PC31DOWNTO2_intermed_5 <= R_D_PC31DOWNTO2_intermed_4;
		R_D_PC31DOWNTO2_intermed_6 <= R_D_PC31DOWNTO2_intermed_5;
		RIN_F_PC31DOWNTO2_intermed_1 <= RIN.F.PC ( 31 DOWNTO 2 );
		IR_ADDR31DOWNTO2_intermed_1 <= IR.ADDR( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_4 <= RIN_E_CTRL_PC31DOWNTO2_intermed_3;
		RIN_E_CTRL_PC31DOWNTO2_intermed_5 <= RIN_E_CTRL_PC31DOWNTO2_intermed_4;
		R_F_PC31DOWNTO2_intermed_1 <= R.F.PC( 31 DOWNTO 2 );
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO2_shadow;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_2;
		VIR_ADDR31DOWNTO2_shadow_intermed_1 <= VIR_ADDR31DOWNTO2_shadow;
		VIR_ADDR31DOWNTO2_shadow_intermed_2 <= VIR_ADDR31DOWNTO2_shadow_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 2 );
		R_M_CTRL_PC31DOWNTO2_intermed_2 <= R_M_CTRL_PC31DOWNTO2_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_3 <= R_M_CTRL_PC31DOWNTO2_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_3 <= RIN_M_CTRL_PC31DOWNTO2_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_4 <= RIN_M_CTRL_PC31DOWNTO2_intermed_3;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_4;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		RIN_A_CTRL_PC31DOWNTO2_intermed_5 <= RIN_A_CTRL_PC31DOWNTO2_intermed_4;
		RIN_A_CTRL_PC31DOWNTO2_intermed_6 <= RIN_A_CTRL_PC31DOWNTO2_intermed_5;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_4 <= R_A_CTRL_PC31DOWNTO2_intermed_3;
		R_A_CTRL_PC31DOWNTO2_intermed_5 <= R_A_CTRL_PC31DOWNTO2_intermed_4;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_3;
		R_X_CTRL_PC31DOWNTO2_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 2 );
		R_X_CTRL_PC31DOWNTO2_intermed_2 <= R_X_CTRL_PC31DOWNTO2_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_5 <= V_D_PC31DOWNTO2_shadow_intermed_4;
		V_D_PC31DOWNTO2_shadow_intermed_6 <= V_D_PC31DOWNTO2_shadow_intermed_5;
		V_D_PC31DOWNTO2_shadow_intermed_7 <= V_D_PC31DOWNTO2_shadow_intermed_6;
		XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_1 <= XC_TRAP_ADDRESS31DOWNTO2_shadow;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_5 <= RIN_D_PC31DOWNTO2_intermed_4;
		RIN_D_PC31DOWNTO2_intermed_6 <= RIN_D_PC31DOWNTO2_intermed_5;
		RIN_D_PC31DOWNTO2_intermed_7 <= RIN_D_PC31DOWNTO2_intermed_6;
		EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_1 <= EX_ADD_RES32DOWNTO332DOWNTO3_shadow;
		V_F_PC31DOWNTO2_shadow_intermed_1 <= V_F_PC31DOWNTO2_shadow;
		RIN_F_PC31DOWNTO2_intermed_1 <= RIN.F.PC( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_2 <= RIN_X_CTRL_PC31DOWNTO2_intermed_1;
		RIN_X_CTRL_PC31DOWNTO2_intermed_3 <= RIN_X_CTRL_PC31DOWNTO2_intermed_2;
		IRIN_ADDR31DOWNTO2_intermed_1 <= IRIN.ADDR( 31 DOWNTO 2 );
		IRIN_ADDR31DOWNTO2_intermed_2 <= IRIN_ADDR31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_3 <= R_E_CTRL_PC31DOWNTO2_intermed_2;
		R_E_CTRL_PC31DOWNTO2_intermed_4 <= R_E_CTRL_PC31DOWNTO2_intermed_3;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_6 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_5;
		EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_1 <= EX_JUMP_ADDRESS31DOWNTO2_shadow;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		R_D_PC31DOWNTO2_intermed_4 <= R_D_PC31DOWNTO2_intermed_3;
		R_D_PC31DOWNTO2_intermed_5 <= R_D_PC31DOWNTO2_intermed_4;
		R_D_PC31DOWNTO2_intermed_6 <= R_D_PC31DOWNTO2_intermed_5;
		IR_ADDR31DOWNTO2_intermed_1 <= IR.ADDR( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_4 <= RIN_E_CTRL_PC31DOWNTO2_intermed_3;
		RIN_E_CTRL_PC31DOWNTO2_intermed_5 <= RIN_E_CTRL_PC31DOWNTO2_intermed_4;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO2_shadow;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_2;
		VIR_ADDR31DOWNTO2_shadow_intermed_1 <= VIR_ADDR31DOWNTO2_shadow;
		VIR_ADDR31DOWNTO2_shadow_intermed_2 <= VIR_ADDR31DOWNTO2_shadow_intermed_1;
		V_X_ANNUL_ALL_shadow_intermed_1 <= V_X_ANNUL_ALL_shadow;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		V_A_MULSTART_shadow_intermed_1 <= V_A_MULSTART_shadow;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_X_ANNUL_ALL_intermed_2 <= RIN_X_ANNUL_ALL_intermed_1;
		R_X_ANNUL_ALL_intermed_1 <= R.X.ANNUL_ALL;
		RIN_A_MULSTART_intermed_1 <= RIN.A.MULSTART;
		V_A_CTRL_ANNUL_shadow_intermed_1 <= V_A_CTRL_ANNUL_shadow;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA ( 0 )( 31 );
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		V_X_DATA0_shadow_intermed_2 <= V_X_DATA0_shadow_intermed_1;
		DE_INST19_shadow_intermed_1 <= DE_INST19_shadow;
		DE_INST19_shadow_intermed_2 <= DE_INST19_shadow_intermed_1;
		RIN_E_OP131_intermed_1 <= RIN.E.OP1( 31 );
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_3 <= V_A_CTRL_INST19_shadow_intermed_2;
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA ( 0 );
		V_E_OP131_shadow_intermed_1 <= V_E_OP131_shadow;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_E_CTRL_INST19_shadow_intermed_1 <= V_E_CTRL_INST19_shadow;
		V_E_OP1_shadow_intermed_1 <= V_E_OP1_shadow;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_2 <= V_X_DATA031_shadow_intermed_1;
		V_E_CTRL_INST19_shadow_intermed_1 <= V_E_CTRL_INST19_shadow;
		V_E_CTRL_INST19_shadow_intermed_2 <= V_E_CTRL_INST19_shadow_intermed_1;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA( 0 )( 31 );
		RIN_X_DATA031_intermed_2 <= RIN_X_DATA031_intermed_1;
		RIN_E_OP1_intermed_1 <= RIN.E.OP1;
		R_E_CTRL_INST19_intermed_1 <= R.E.CTRL.INST( 19 );
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		DCO_DATA031_intermed_1 <= DCO.DATA ( 0 )( 31 );
		R_X_DATA031_intermed_1 <= R.X.DATA( 0 )( 31 );
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST ( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		R_X_DATA0_intermed_1 <= R.X.DATA( 0 );
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST( 19 );
		R_A_CTRL_INST19_intermed_2 <= R_A_CTRL_INST19_intermed_1;
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST ( 19 );
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		RIN_A_CTRL_INST19_intermed_3 <= RIN_A_CTRL_INST19_intermed_2;
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST ( 19 );
		DCO_DATA0_intermed_1 <= DCO.DATA ( 0 );
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA( 0 );
		RIN_X_DATA0_intermed_2 <= RIN_X_DATA0_intermed_1;
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST( 19 );
		RIN_E_CTRL_INST19_intermed_2 <= RIN_E_CTRL_INST19_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA ( 0 )( 31 );
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		V_X_DATA0_shadow_intermed_2 <= V_X_DATA0_shadow_intermed_1;
		DE_INST19_shadow_intermed_1 <= DE_INST19_shadow;
		DE_INST19_shadow_intermed_2 <= DE_INST19_shadow_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_3 <= V_A_CTRL_INST19_shadow_intermed_2;
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA ( 0 );
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_E_CTRL_INST19_shadow_intermed_1 <= V_E_CTRL_INST19_shadow;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_2 <= V_X_DATA031_shadow_intermed_1;
		V_E_OP2_shadow_intermed_1 <= V_E_OP2_shadow;
		RIN_E_OP2_intermed_1 <= RIN.E.OP2;
		V_E_CTRL_INST19_shadow_intermed_1 <= V_E_CTRL_INST19_shadow;
		V_E_CTRL_INST19_shadow_intermed_2 <= V_E_CTRL_INST19_shadow_intermed_1;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA( 0 )( 31 );
		RIN_X_DATA031_intermed_2 <= RIN_X_DATA031_intermed_1;
		R_E_CTRL_INST19_intermed_1 <= R.E.CTRL.INST( 19 );
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		DCO_DATA031_intermed_1 <= DCO.DATA ( 0 )( 31 );
		R_X_DATA031_intermed_1 <= R.X.DATA( 0 )( 31 );
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST ( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		R_X_DATA0_intermed_1 <= R.X.DATA( 0 );
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST( 19 );
		R_A_CTRL_INST19_intermed_2 <= R_A_CTRL_INST19_intermed_1;
		RIN_E_OP231_intermed_1 <= RIN.E.OP2( 31 );
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST ( 19 );
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		RIN_A_CTRL_INST19_intermed_3 <= RIN_A_CTRL_INST19_intermed_2;
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST ( 19 );
		V_E_OP231_shadow_intermed_1 <= V_E_OP231_shadow;
		DCO_DATA0_intermed_1 <= DCO.DATA ( 0 );
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA( 0 );
		RIN_X_DATA0_intermed_2 <= RIN_X_DATA0_intermed_1;
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST( 19 );
		RIN_E_CTRL_INST19_intermed_2 <= RIN_E_CTRL_INST19_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		V_A_CTRL_INST24_shadow_intermed_1 <= V_A_CTRL_INST24_shadow;
		V_A_CTRL_INST24_shadow_intermed_2 <= V_A_CTRL_INST24_shadow_intermed_1;
		V_A_CTRL_INST24_shadow_intermed_3 <= V_A_CTRL_INST24_shadow_intermed_2;
		V_E_CTRL_INST24_shadow_intermed_1 <= V_E_CTRL_INST24_shadow;
		V_E_CTRL_INST24_shadow_intermed_2 <= V_E_CTRL_INST24_shadow_intermed_1;
		DE_INST24_shadow_intermed_1 <= DE_INST24_shadow;
		DE_INST24_shadow_intermed_2 <= DE_INST24_shadow_intermed_1;
		DE_INST24_shadow_intermed_3 <= DE_INST24_shadow_intermed_2;
		V_E_CTRL_INST24_shadow_intermed_1 <= V_E_CTRL_INST24_shadow;
		R_A_CTRL_INST24_intermed_1 <= R.A.CTRL.INST( 24 );
		R_A_CTRL_INST24_intermed_2 <= R_A_CTRL_INST24_intermed_1;
		RIN_A_CTRL_INST24_intermed_1 <= RIN.A.CTRL.INST ( 24 );
		RIN_A_CTRL_INST24_intermed_2 <= RIN_A_CTRL_INST24_intermed_1;
		V_A_CTRL_INST24_shadow_intermed_1 <= V_A_CTRL_INST24_shadow;
		V_A_CTRL_INST24_shadow_intermed_2 <= V_A_CTRL_INST24_shadow_intermed_1;
		RIN_A_CTRL_INST24_intermed_1 <= RIN.A.CTRL.INST( 24 );
		RIN_A_CTRL_INST24_intermed_2 <= RIN_A_CTRL_INST24_intermed_1;
		RIN_A_CTRL_INST24_intermed_3 <= RIN_A_CTRL_INST24_intermed_2;
		RIN_E_CTRL_INST24_intermed_1 <= RIN.E.CTRL.INST( 24 );
		RIN_E_CTRL_INST24_intermed_2 <= RIN_E_CTRL_INST24_intermed_1;
		R_E_CTRL_INST24_intermed_1 <= R.E.CTRL.INST( 24 );
		R_E_CTRL_INST24_intermed_2 <= R_E_CTRL_INST24_intermed_1;
		R_A_CTRL_INST24_intermed_1 <= R.A.CTRL.INST ( 24 );
		RIN_E_CTRL_INST24_intermed_1 <= RIN.E.CTRL.INST ( 24 );
		V_X_ANNUL_ALL_shadow_intermed_1 <= V_X_ANNUL_ALL_shadow;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_A_DIVSTART_intermed_1 <= RIN.A.DIVSTART;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_X_ANNUL_ALL_intermed_2 <= RIN_X_ANNUL_ALL_intermed_1;
		R_X_ANNUL_ALL_intermed_1 <= R.X.ANNUL_ALL;
		V_A_DIVSTART_shadow_intermed_1 <= V_A_DIVSTART_shadow;
		V_A_CTRL_ANNUL_shadow_intermed_1 <= V_A_CTRL_ANNUL_shadow;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA ( 0 )( 31 );
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		V_X_DATA0_shadow_intermed_2 <= V_X_DATA0_shadow_intermed_1;
		DE_INST19_shadow_intermed_1 <= DE_INST19_shadow;
		DE_INST19_shadow_intermed_2 <= DE_INST19_shadow_intermed_1;
		RIN_E_OP131_intermed_1 <= RIN.E.OP1( 31 );
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_3 <= V_A_CTRL_INST19_shadow_intermed_2;
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA ( 0 );
		V_E_OP131_shadow_intermed_1 <= V_E_OP131_shadow;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_E_CTRL_INST19_shadow_intermed_1 <= V_E_CTRL_INST19_shadow;
		V_E_OP1_shadow_intermed_1 <= V_E_OP1_shadow;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_2 <= V_X_DATA031_shadow_intermed_1;
		V_E_CTRL_INST19_shadow_intermed_1 <= V_E_CTRL_INST19_shadow;
		V_E_CTRL_INST19_shadow_intermed_2 <= V_E_CTRL_INST19_shadow_intermed_1;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA( 0 )( 31 );
		RIN_X_DATA031_intermed_2 <= RIN_X_DATA031_intermed_1;
		RIN_E_OP1_intermed_1 <= RIN.E.OP1;
		R_E_CTRL_INST19_intermed_1 <= R.E.CTRL.INST( 19 );
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		DCO_DATA031_intermed_1 <= DCO.DATA ( 0 )( 31 );
		R_X_DATA031_intermed_1 <= R.X.DATA( 0 )( 31 );
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST ( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		R_X_DATA0_intermed_1 <= R.X.DATA( 0 );
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST( 19 );
		R_A_CTRL_INST19_intermed_2 <= R_A_CTRL_INST19_intermed_1;
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST ( 19 );
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		RIN_A_CTRL_INST19_intermed_3 <= RIN_A_CTRL_INST19_intermed_2;
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST ( 19 );
		DCO_DATA0_intermed_1 <= DCO.DATA ( 0 );
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA( 0 );
		RIN_X_DATA0_intermed_2 <= RIN_X_DATA0_intermed_1;
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST( 19 );
		RIN_E_CTRL_INST19_intermed_2 <= RIN_E_CTRL_INST19_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA ( 0 )( 31 );
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		V_X_DATA0_shadow_intermed_2 <= V_X_DATA0_shadow_intermed_1;
		DE_INST19_shadow_intermed_1 <= DE_INST19_shadow;
		DE_INST19_shadow_intermed_2 <= DE_INST19_shadow_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_3 <= V_A_CTRL_INST19_shadow_intermed_2;
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA ( 0 );
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_E_CTRL_INST19_shadow_intermed_1 <= V_E_CTRL_INST19_shadow;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_2 <= V_X_DATA031_shadow_intermed_1;
		V_E_OP2_shadow_intermed_1 <= V_E_OP2_shadow;
		RIN_E_OP2_intermed_1 <= RIN.E.OP2;
		V_E_CTRL_INST19_shadow_intermed_1 <= V_E_CTRL_INST19_shadow;
		V_E_CTRL_INST19_shadow_intermed_2 <= V_E_CTRL_INST19_shadow_intermed_1;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA( 0 )( 31 );
		RIN_X_DATA031_intermed_2 <= RIN_X_DATA031_intermed_1;
		R_E_CTRL_INST19_intermed_1 <= R.E.CTRL.INST( 19 );
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		DCO_DATA031_intermed_1 <= DCO.DATA ( 0 )( 31 );
		R_X_DATA031_intermed_1 <= R.X.DATA( 0 )( 31 );
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST ( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		R_X_DATA0_intermed_1 <= R.X.DATA( 0 );
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST( 19 );
		R_A_CTRL_INST19_intermed_2 <= R_A_CTRL_INST19_intermed_1;
		RIN_E_OP231_intermed_1 <= RIN.E.OP2( 31 );
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST ( 19 );
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		RIN_A_CTRL_INST19_intermed_3 <= RIN_A_CTRL_INST19_intermed_2;
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST ( 19 );
		V_E_OP231_shadow_intermed_1 <= V_E_OP231_shadow;
		DCO_DATA0_intermed_1 <= DCO.DATA ( 0 );
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA( 0 );
		RIN_X_DATA0_intermed_2 <= RIN_X_DATA0_intermed_1;
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST( 19 );
		RIN_E_CTRL_INST19_intermed_2 <= RIN_E_CTRL_INST19_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		DE_INST19_shadow_intermed_1 <= DE_INST19_shadow;
		DE_INST19_shadow_intermed_2 <= DE_INST19_shadow_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST ( 19 );
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST( 19 );
		R_A_CTRL_INST19_intermed_2 <= R_A_CTRL_INST19_intermed_1;
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		DE_INST19_shadow_intermed_1 <= DE_INST19_shadow;
		RIN_M_Y31_intermed_1 <= RIN.M.Y ( 31 );
		RIN_M_Y_intermed_1 <= RIN.M.Y;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		V_E_CTRL_INST19_shadow_intermed_1 <= V_E_CTRL_INST19_shadow;
		V_M_Y31_shadow_intermed_1 <= V_M_Y31_shadow;
		V_M_Y31_shadow_intermed_2 <= V_M_Y31_shadow_intermed_1;
		V_M_Y_shadow_intermed_1 <= V_M_Y_shadow;
		V_E_CTRL_INST19_shadow_intermed_1 <= V_E_CTRL_INST19_shadow;
		V_E_CTRL_INST19_shadow_intermed_2 <= V_E_CTRL_INST19_shadow_intermed_1;
		R_E_CTRL_INST19_intermed_1 <= R.E.CTRL.INST( 19 );
		V_M_Y31_shadow_intermed_1 <= V_M_Y31_shadow;
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST ( 19 );
		RIN_M_Y31_intermed_1 <= RIN.M.Y( 31 );
		RIN_M_Y31_intermed_2 <= RIN_M_Y31_intermed_1;
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST( 19 );
		R_M_Y31_intermed_1 <= R.M.Y( 31 );
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST ( 19 );
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST( 19 );
		RIN_E_CTRL_INST19_intermed_2 <= RIN_E_CTRL_INST19_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		RIN_M_Y31_intermed_1 <= RIN.M.Y ( 31 );
		V_M_Y31_shadow_intermed_1 <= V_M_Y31_shadow;
		V_M_Y31_shadow_intermed_2 <= V_M_Y31_shadow_intermed_1;
		V_M_Y31_shadow_intermed_1 <= V_M_Y31_shadow;
		RIN_M_Y31_intermed_1 <= RIN.M.Y( 31 );
		RIN_M_Y31_intermed_2 <= RIN_M_Y31_intermed_1;
		R_M_Y31_intermed_1 <= R.M.Y( 31 );
		R_M_Y31_intermed_2 <= R_M_Y31_intermed_1;
		VDSU_CRDY2_shadow_intermed_1 <= VDSU_CRDY2_shadow;
		VDSU_CRDY2_shadow_intermed_2 <= VDSU_CRDY2_shadow_intermed_1;
		DSUIN_CRDY2_intermed_1 <= DSUIN.CRDY ( 2 );
		VDSU_CRDY2_shadow_intermed_1 <= VDSU_CRDY2_shadow;
		DSUIN_CRDY2_intermed_1 <= DSUIN.CRDY( 2 );
		DSUIN_CRDY2_intermed_2 <= DSUIN_CRDY2_intermed_1;
		DSUR_CRDY2_intermed_1 <= DSUR.CRDY( 2 );
		DSUR_CRDY2_intermed_2 <= DSUR_CRDY2_intermed_1;
		VP_ERROR_shadow_intermed_1 <= VP_ERROR_shadow;
		VP_ERROR_shadow_intermed_2 <= VP_ERROR_shadow_intermed_1;
		RIN_X_NERROR_intermed_1 <= RIN.X.NERROR;
		RPIN_ERROR_intermed_1 <= RPIN.ERROR;
		RPIN_ERROR_intermed_2 <= RPIN_ERROR_intermed_1;
		V_X_NERROR_shadow_intermed_1 <= V_X_NERROR_shadow;
		RP_ERROR_intermed_1 <= RP.ERROR;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC ( 31 DOWNTO 2 );
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC ( 31 DOWNTO 2 );
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC ( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC ( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 2 );
		R_M_CTRL_PC31DOWNTO2_intermed_2 <= R_M_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC ( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC ( 31 DOWNTO 2 );
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_5 <= V_D_PC31DOWNTO2_shadow_intermed_4;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_5 <= RIN_D_PC31DOWNTO2_intermed_4;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC ( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC ( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC ( 31 DOWNTO 2 );
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		R_D_PC31DOWNTO2_intermed_4 <= R_D_PC31DOWNTO2_intermed_3;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_X_RESULT6DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO0_shadow;
		RIN_X_RESULT6DOWNTO0_intermed_1 <= RIN.X.RESULT( 6 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO0_intermed_2 <= RIN_X_RESULT6DOWNTO0_intermed_1;
		R_X_RESULT6DOWNTO0_intermed_1 <= R.X.RESULT( 6 DOWNTO 0 );
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		R_X_DATA0_intermed_1 <= R.X.DATA( 0 );
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA( 0 );
		RIN_X_DATA0_intermed_2 <= RIN_X_DATA0_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC ( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC ( 31 DOWNTO 2 );
		R_X_CTRL_PC31DOWNTO2_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 2 );
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_5 <= V_D_PC31DOWNTO2_shadow_intermed_4;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_5 <= RIN_D_PC31DOWNTO2_intermed_4;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC ( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC ( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC ( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_2 <= RIN_X_CTRL_PC31DOWNTO2_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		R_D_PC31DOWNTO2_intermed_4 <= R_D_PC31DOWNTO2_intermed_3;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO2_shadow;
		V_X_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_X_CTRL_TT3DOWNTO0_shadow;
		V_X_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_X_CTRL_TT3DOWNTO0_shadow_intermed_1;
		R_M_CTRL_TT3DOWNTO0_intermed_1 <= R.M.CTRL.TT( 3 DOWNTO 0 );
		R_M_CTRL_TT3DOWNTO0_intermed_2 <= R_M_CTRL_TT3DOWNTO0_intermed_1;
		V_M_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_M_CTRL_TT3DOWNTO0_shadow;
		V_M_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_M_CTRL_TT3DOWNTO0_shadow_intermed_1;
		V_M_CTRL_TT3DOWNTO0_shadow_intermed_3 <= V_M_CTRL_TT3DOWNTO0_shadow_intermed_2;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_3 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2;
		R_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= R.X.RESULT( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		R_X_RESULT6DOWNTO03DOWNTO0_intermed_2 <= R_X_RESULT6DOWNTO03DOWNTO0_intermed_1;
		R_A_CTRL_TT3DOWNTO0_intermed_1 <= R.A.CTRL.TT( 3 DOWNTO 0 );
		R_A_CTRL_TT3DOWNTO0_intermed_2 <= R_A_CTRL_TT3DOWNTO0_intermed_1;
		R_A_CTRL_TT3DOWNTO0_intermed_3 <= R_A_CTRL_TT3DOWNTO0_intermed_2;
		R_A_CTRL_TT3DOWNTO0_intermed_4 <= R_A_CTRL_TT3DOWNTO0_intermed_3;
		RIN_A_CTRL_TT3DOWNTO0_intermed_1 <= RIN.A.CTRL.TT( 3 DOWNTO 0 );
		RIN_A_CTRL_TT3DOWNTO0_intermed_2 <= RIN_A_CTRL_TT3DOWNTO0_intermed_1;
		RIN_A_CTRL_TT3DOWNTO0_intermed_3 <= RIN_A_CTRL_TT3DOWNTO0_intermed_2;
		RIN_A_CTRL_TT3DOWNTO0_intermed_4 <= RIN_A_CTRL_TT3DOWNTO0_intermed_3;
		RIN_A_CTRL_TT3DOWNTO0_intermed_5 <= RIN_A_CTRL_TT3DOWNTO0_intermed_4;
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= RIN.X.RESULT( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2 <= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1;
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_3 <= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_A_CTRL_TT3DOWNTO0_shadow;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_1;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_3 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_2;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_4 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_3;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_5 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_4;
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= RIN.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2 <= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1;
		R_W_S_TT3DOWNTO0_intermed_1 <= R.W.S.TT( 3 DOWNTO 0 );
		R_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= R.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		R_E_CTRL_TT3DOWNTO0_intermed_1 <= R.E.CTRL.TT( 3 DOWNTO 0 );
		R_E_CTRL_TT3DOWNTO0_intermed_2 <= R_E_CTRL_TT3DOWNTO0_intermed_1;
		R_E_CTRL_TT3DOWNTO0_intermed_3 <= R_E_CTRL_TT3DOWNTO0_intermed_2;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1;
		RIN_W_S_TT3DOWNTO0_intermed_1 <= RIN.W.S.TT( 3 DOWNTO 0 );
		RIN_W_S_TT3DOWNTO0_intermed_2 <= RIN_W_S_TT3DOWNTO0_intermed_1;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_E_CTRL_TT3DOWNTO0_shadow;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_E_CTRL_TT3DOWNTO0_shadow_intermed_1;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_3 <= V_E_CTRL_TT3DOWNTO0_shadow_intermed_2;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_4 <= V_E_CTRL_TT3DOWNTO0_shadow_intermed_3;
		RIN_M_CTRL_TT3DOWNTO0_intermed_1 <= RIN.M.CTRL.TT( 3 DOWNTO 0 );
		RIN_M_CTRL_TT3DOWNTO0_intermed_2 <= RIN_M_CTRL_TT3DOWNTO0_intermed_1;
		RIN_M_CTRL_TT3DOWNTO0_intermed_3 <= RIN_M_CTRL_TT3DOWNTO0_intermed_2;
		RIN_X_CTRL_TT3DOWNTO0_intermed_1 <= RIN.X.CTRL.TT( 3 DOWNTO 0 );
		RIN_X_CTRL_TT3DOWNTO0_intermed_2 <= RIN_X_CTRL_TT3DOWNTO0_intermed_1;
		V_W_S_TT3DOWNTO0_shadow_intermed_1 <= V_W_S_TT3DOWNTO0_shadow;
		R_X_CTRL_TT3DOWNTO0_intermed_1 <= R.X.CTRL.TT( 3 DOWNTO 0 );
		RIN_E_CTRL_TT3DOWNTO0_intermed_1 <= RIN.E.CTRL.TT( 3 DOWNTO 0 );
		RIN_E_CTRL_TT3DOWNTO0_intermed_2 <= RIN_E_CTRL_TT3DOWNTO0_intermed_1;
		RIN_E_CTRL_TT3DOWNTO0_intermed_3 <= RIN_E_CTRL_TT3DOWNTO0_intermed_2;
		RIN_E_CTRL_TT3DOWNTO0_intermed_4 <= RIN_E_CTRL_TT3DOWNTO0_intermed_3;
		XC_VECTT3DOWNTO0_shadow_intermed_1 <= XC_VECTT3DOWNTO0_shadow;
		V_M_RESULT1DOWNTO0_shadow_intermed_1 <= V_M_RESULT1DOWNTO0_shadow;
		RIN_M_RESULT1DOWNTO0_intermed_1 <= RIN.M.RESULT( 1 DOWNTO 0 );
		RIN_M_RESULT1DOWNTO0_intermed_2 <= RIN_M_RESULT1DOWNTO0_intermed_1;
		R_M_RESULT1DOWNTO0_intermed_1 <= R.M.RESULT( 1 DOWNTO 0 );
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA ( 0 )( 31 );
		RIN_X_DATA031_intermed_2 <= RIN_X_DATA031_intermed_1;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA( 0 )( 31 );
		RIN_X_DATA031_intermed_2 <= RIN_X_DATA031_intermed_1;
		DCO_DATA031_intermed_1 <= DCO.DATA ( 0 )( 31 );
		R_X_DATA031_intermed_1 <= R.X.DATA( 0 )( 31 );
		R_X_DATA031_intermed_1 <= R.X.DATA ( 0 )( 31 );
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA( 0 )( 31 );
		RIN_X_DATA031_intermed_2 <= RIN_X_DATA031_intermed_1;
		R_X_DATA031_intermed_1 <= R.X.DATA( 0 )( 31 );
		DE_INST19_shadow_intermed_1 <= DE_INST19_shadow;
		DE_INST19_shadow_intermed_2 <= DE_INST19_shadow_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		V_E_CTRL_INST19_shadow_intermed_1 <= V_E_CTRL_INST19_shadow;
		R_E_CTRL_INST19_intermed_1 <= R.E.CTRL.INST( 19 );
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST ( 19 );
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST( 19 );
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST( 19 );
		RIN_E_CTRL_INST19_intermed_2 <= RIN_E_CTRL_INST19_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST20_shadow_intermed_1 <= V_A_CTRL_INST20_shadow;
		RIN_A_CTRL_INST20_intermed_1 <= RIN.A.CTRL.INST ( 20 );
		R_E_CTRL_INST20_intermed_1 <= R.E.CTRL.INST( 20 );
		RIN_A_CTRL_INST20_intermed_1 <= RIN.A.CTRL.INST( 20 );
		RIN_A_CTRL_INST20_intermed_2 <= RIN_A_CTRL_INST20_intermed_1;
		V_E_CTRL_INST20_shadow_intermed_1 <= V_E_CTRL_INST20_shadow;
		DE_INST20_shadow_intermed_1 <= DE_INST20_shadow;
		DE_INST20_shadow_intermed_2 <= DE_INST20_shadow_intermed_1;
		V_A_CTRL_INST20_shadow_intermed_1 <= V_A_CTRL_INST20_shadow;
		V_A_CTRL_INST20_shadow_intermed_2 <= V_A_CTRL_INST20_shadow_intermed_1;
		RIN_E_CTRL_INST20_intermed_1 <= RIN.E.CTRL.INST( 20 );
		RIN_E_CTRL_INST20_intermed_2 <= RIN_E_CTRL_INST20_intermed_1;
		R_A_CTRL_INST20_intermed_1 <= R.A.CTRL.INST( 20 );
		RIN_X_DATA00_intermed_1 <= RIN.X.DATA ( 0 )( 0 );
		RIN_X_DATA00_intermed_2 <= RIN_X_DATA00_intermed_1;
		DCO_DATA00_intermed_1 <= DCO.DATA ( 0 )( 0 );
		V_X_DATA00_shadow_intermed_1 <= V_X_DATA00_shadow;
		V_X_DATA00_shadow_intermed_1 <= V_X_DATA00_shadow;
		R_X_DATA00_intermed_1 <= R.X.DATA ( 0 )( 0 );
		RIN_X_DATA00_intermed_1 <= RIN.X.DATA( 0 )( 0 );
		RIN_X_DATA00_intermed_2 <= RIN_X_DATA00_intermed_1;
		R_X_DATA00_intermed_1 <= R.X.DATA( 0 )( 0 );
		V_X_DATA00_shadow_intermed_1 <= V_X_DATA00_shadow;
		RIN_X_DATA00_intermed_1 <= RIN.X.DATA( 0 )( 0 );
		RIN_X_DATA00_intermed_2 <= RIN_X_DATA00_intermed_1;
		R_X_DATA00_intermed_1 <= R.X.DATA( 0 )( 0 );
		V_X_DATA04DOWNTO0_shadow_intermed_1 <= V_X_DATA04DOWNTO0_shadow;
		R_X_DATA04DOWNTO0_intermed_1 <= R.X.DATA( 0 )( 4 DOWNTO 0 );
		R_X_DATA04DOWNTO0_intermed_1 <= R.X.DATA ( 0 )( 4 DOWNTO 0 );
		DCO_DATA04DOWNTO0_intermed_1 <= DCO.DATA ( 0 )( 4 DOWNTO 0 );
		RIN_X_DATA04DOWNTO0_intermed_1 <= RIN.X.DATA ( 0 )( 4 DOWNTO 0 );
		RIN_X_DATA04DOWNTO0_intermed_2 <= RIN_X_DATA04DOWNTO0_intermed_1;
		RIN_X_DATA04DOWNTO0_intermed_1 <= RIN.X.DATA( 0 )( 4 DOWNTO 0 );
		RIN_X_DATA04DOWNTO0_intermed_2 <= RIN_X_DATA04DOWNTO0_intermed_1;
		V_X_DATA04DOWNTO0_shadow_intermed_1 <= V_X_DATA04DOWNTO0_shadow;
		V_X_DATA04DOWNTO0_shadow_intermed_1 <= V_X_DATA04DOWNTO0_shadow;
		R_X_DATA04DOWNTO0_intermed_1 <= R.X.DATA( 0 )( 4 DOWNTO 0 );
		RIN_X_DATA04DOWNTO0_intermed_1 <= RIN.X.DATA( 0 )( 4 DOWNTO 0 );
		RIN_X_DATA04DOWNTO0_intermed_2 <= RIN_X_DATA04DOWNTO0_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 2 );
		R_M_CTRL_PC31DOWNTO2_intermed_2 <= R_M_CTRL_PC31DOWNTO2_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_3 <= R_M_CTRL_PC31DOWNTO2_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_3 <= RIN_M_CTRL_PC31DOWNTO2_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_4 <= RIN_M_CTRL_PC31DOWNTO2_intermed_3;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_4;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		RIN_A_CTRL_PC31DOWNTO2_intermed_5 <= RIN_A_CTRL_PC31DOWNTO2_intermed_4;
		RIN_A_CTRL_PC31DOWNTO2_intermed_6 <= RIN_A_CTRL_PC31DOWNTO2_intermed_5;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_4 <= R_A_CTRL_PC31DOWNTO2_intermed_3;
		R_A_CTRL_PC31DOWNTO2_intermed_5 <= R_A_CTRL_PC31DOWNTO2_intermed_4;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_3;
		R_X_CTRL_PC31DOWNTO2_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 2 );
		R_X_CTRL_PC31DOWNTO2_intermed_2 <= R_X_CTRL_PC31DOWNTO2_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_5 <= V_D_PC31DOWNTO2_shadow_intermed_4;
		V_D_PC31DOWNTO2_shadow_intermed_6 <= V_D_PC31DOWNTO2_shadow_intermed_5;
		V_D_PC31DOWNTO2_shadow_intermed_7 <= V_D_PC31DOWNTO2_shadow_intermed_6;
		XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_1 <= XC_TRAP_ADDRESS31DOWNTO2_shadow;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_5 <= RIN_D_PC31DOWNTO2_intermed_4;
		RIN_D_PC31DOWNTO2_intermed_6 <= RIN_D_PC31DOWNTO2_intermed_5;
		RIN_D_PC31DOWNTO2_intermed_7 <= RIN_D_PC31DOWNTO2_intermed_6;
		EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_1 <= EX_ADD_RES32DOWNTO332DOWNTO3_shadow;
		V_F_PC31DOWNTO2_shadow_intermed_1 <= V_F_PC31DOWNTO2_shadow;
		RIN_F_PC31DOWNTO2_intermed_1 <= RIN.F.PC( 31 DOWNTO 2 );
		RIN_F_PC31DOWNTO2_intermed_2 <= RIN_F_PC31DOWNTO2_intermed_1;
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_2 <= RIN_X_CTRL_PC31DOWNTO2_intermed_1;
		RIN_X_CTRL_PC31DOWNTO2_intermed_3 <= RIN_X_CTRL_PC31DOWNTO2_intermed_2;
		IRIN_ADDR31DOWNTO2_intermed_1 <= IRIN.ADDR( 31 DOWNTO 2 );
		IRIN_ADDR31DOWNTO2_intermed_2 <= IRIN_ADDR31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_3 <= R_E_CTRL_PC31DOWNTO2_intermed_2;
		R_E_CTRL_PC31DOWNTO2_intermed_4 <= R_E_CTRL_PC31DOWNTO2_intermed_3;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_6 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_5;
		EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_1 <= EX_JUMP_ADDRESS31DOWNTO2_shadow;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		R_D_PC31DOWNTO2_intermed_4 <= R_D_PC31DOWNTO2_intermed_3;
		R_D_PC31DOWNTO2_intermed_5 <= R_D_PC31DOWNTO2_intermed_4;
		R_D_PC31DOWNTO2_intermed_6 <= R_D_PC31DOWNTO2_intermed_5;
		IR_ADDR31DOWNTO2_intermed_1 <= IR.ADDR( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_4 <= RIN_E_CTRL_PC31DOWNTO2_intermed_3;
		RIN_E_CTRL_PC31DOWNTO2_intermed_5 <= RIN_E_CTRL_PC31DOWNTO2_intermed_4;
		R_F_PC31DOWNTO2_intermed_1 <= R.F.PC( 31 DOWNTO 2 );
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO2_shadow;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_2;
		VIR_ADDR31DOWNTO2_shadow_intermed_1 <= VIR_ADDR31DOWNTO2_shadow;
		VIR_ADDR31DOWNTO2_shadow_intermed_2 <= VIR_ADDR31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		V_A_CTRL_INST24_shadow_intermed_1 <= V_A_CTRL_INST24_shadow;
		V_A_CTRL_INST24_shadow_intermed_2 <= V_A_CTRL_INST24_shadow_intermed_1;
		V_E_CTRL_INST24_shadow_intermed_1 <= V_E_CTRL_INST24_shadow;
		DE_INST24_shadow_intermed_1 <= DE_INST24_shadow;
		DE_INST24_shadow_intermed_2 <= DE_INST24_shadow_intermed_1;
		R_A_CTRL_INST24_intermed_1 <= R.A.CTRL.INST( 24 );
		RIN_A_CTRL_INST24_intermed_1 <= RIN.A.CTRL.INST ( 24 );
		V_A_CTRL_INST24_shadow_intermed_1 <= V_A_CTRL_INST24_shadow;
		RIN_A_CTRL_INST24_intermed_1 <= RIN.A.CTRL.INST( 24 );
		RIN_A_CTRL_INST24_intermed_2 <= RIN_A_CTRL_INST24_intermed_1;
		RIN_E_CTRL_INST24_intermed_1 <= RIN.E.CTRL.INST( 24 );
		RIN_E_CTRL_INST24_intermed_2 <= RIN_E_CTRL_INST24_intermed_1;
		R_E_CTRL_INST24_intermed_1 <= R.E.CTRL.INST( 24 );
		DE_INST19_shadow_intermed_1 <= DE_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST( 19 );
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		V_M_Y31_shadow_intermed_1 <= V_M_Y31_shadow;
		RIN_M_Y31_intermed_1 <= RIN.M.Y( 31 );
		RIN_M_Y31_intermed_2 <= RIN_M_Y31_intermed_1;
		R_M_Y31_intermed_1 <= R.M.Y( 31 );
		VDSU_CRDY2_shadow_intermed_1 <= VDSU_CRDY2_shadow;
		DSUIN_CRDY2_intermed_1 <= DSUIN.CRDY( 2 );
		DSUIN_CRDY2_intermed_2 <= DSUIN_CRDY2_intermed_1;
		DSUR_CRDY2_intermed_1 <= DSUR.CRDY( 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC ( 31 DOWNTO 2 );
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC ( 31 DOWNTO 2 );
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC ( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC ( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_X_DATA1_shadow_intermed_1 <= V_X_DATA1_shadow;
		DCO_DATA1_intermed_1 <= DCO.DATA ( 1 );
		V_X_DATA1_shadow_intermed_1 <= V_X_DATA1_shadow;
		V_X_DATA1_shadow_intermed_2 <= V_X_DATA1_shadow_intermed_1;
		RIN_X_DATA1_intermed_1 <= RIN.X.DATA ( 1 );
		R_X_DATA1_intermed_1 <= R.X.DATA( 1 );
		R_X_DATA1_intermed_2 <= R_X_DATA1_intermed_1;
		RIN_X_DATA1_intermed_1 <= RIN.X.DATA( 1 );
		RIN_X_DATA1_intermed_2 <= RIN_X_DATA1_intermed_1;
		EX_JUMP_ADDRESS31DOWNTO12_shadow_intermed_1 <= EX_JUMP_ADDRESS31DOWNTO12_shadow;
		EX_JUMP_ADDRESS31DOWNTO12_shadow_intermed_2 <= EX_JUMP_ADDRESS31DOWNTO12_shadow_intermed_1;
		RIN_F_PC31DOWNTO12_intermed_1 <= RIN.F.PC ( 31 DOWNTO 12 );
		RIN_A_CTRL_PC31DOWNTO12_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 12 );
		RIN_A_CTRL_PC31DOWNTO12_intermed_2 <= RIN_A_CTRL_PC31DOWNTO12_intermed_1;
		RIN_A_CTRL_PC31DOWNTO12_intermed_3 <= RIN_A_CTRL_PC31DOWNTO12_intermed_2;
		RIN_A_CTRL_PC31DOWNTO12_intermed_4 <= RIN_A_CTRL_PC31DOWNTO12_intermed_3;
		RIN_A_CTRL_PC31DOWNTO12_intermed_5 <= RIN_A_CTRL_PC31DOWNTO12_intermed_4;
		RIN_A_CTRL_PC31DOWNTO12_intermed_6 <= RIN_A_CTRL_PC31DOWNTO12_intermed_5;
		RIN_A_CTRL_PC31DOWNTO12_intermed_7 <= RIN_A_CTRL_PC31DOWNTO12_intermed_6;
		RIN_E_CTRL_PC31DOWNTO12_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 12 );
		RIN_E_CTRL_PC31DOWNTO12_intermed_2 <= RIN_E_CTRL_PC31DOWNTO12_intermed_1;
		RIN_E_CTRL_PC31DOWNTO12_intermed_3 <= RIN_E_CTRL_PC31DOWNTO12_intermed_2;
		RIN_E_CTRL_PC31DOWNTO12_intermed_4 <= RIN_E_CTRL_PC31DOWNTO12_intermed_3;
		RIN_E_CTRL_PC31DOWNTO12_intermed_5 <= RIN_E_CTRL_PC31DOWNTO12_intermed_4;
		RIN_E_CTRL_PC31DOWNTO12_intermed_6 <= RIN_E_CTRL_PC31DOWNTO12_intermed_5;
		V_F_PC31DOWNTO12_shadow_intermed_1 <= V_F_PC31DOWNTO12_shadow;
		V_F_PC31DOWNTO12_shadow_intermed_2 <= V_F_PC31DOWNTO12_shadow_intermed_1;
		R_M_CTRL_PC31DOWNTO12_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 12 );
		R_M_CTRL_PC31DOWNTO12_intermed_2 <= R_M_CTRL_PC31DOWNTO12_intermed_1;
		R_M_CTRL_PC31DOWNTO12_intermed_3 <= R_M_CTRL_PC31DOWNTO12_intermed_2;
		R_M_CTRL_PC31DOWNTO12_intermed_4 <= R_M_CTRL_PC31DOWNTO12_intermed_3;
		IRIN_ADDR31DOWNTO12_intermed_1 <= IRIN.ADDR( 31 DOWNTO 12 );
		IRIN_ADDR31DOWNTO12_intermed_2 <= IRIN_ADDR31DOWNTO12_intermed_1;
		IRIN_ADDR31DOWNTO12_intermed_3 <= IRIN_ADDR31DOWNTO12_intermed_2;
		V_X_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO12_shadow;
		V_X_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_X_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_X_CTRL_PC31DOWNTO12_shadow_intermed_4 <= V_X_CTRL_PC31DOWNTO12_shadow_intermed_3;
		EX_ADD_RES32DOWNTO332DOWNTO13_shadow_intermed_1 <= EX_ADD_RES32DOWNTO332DOWNTO13_shadow;
		EX_ADD_RES32DOWNTO332DOWNTO13_shadow_intermed_2 <= EX_ADD_RES32DOWNTO332DOWNTO13_shadow_intermed_1;
		XC_TRAP_ADDRESS31DOWNTO12_shadow_intermed_1 <= XC_TRAP_ADDRESS31DOWNTO12_shadow;
		XC_TRAP_ADDRESS31DOWNTO12_shadow_intermed_2 <= XC_TRAP_ADDRESS31DOWNTO12_shadow_intermed_1;
		R_F_PC31DOWNTO12_intermed_1 <= R.F.PC( 31 DOWNTO 12 );
		R_F_PC31DOWNTO12_intermed_2 <= R_F_PC31DOWNTO12_intermed_1;
		RIN_M_CTRL_PC31DOWNTO12_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 12 );
		RIN_M_CTRL_PC31DOWNTO12_intermed_2 <= RIN_M_CTRL_PC31DOWNTO12_intermed_1;
		RIN_M_CTRL_PC31DOWNTO12_intermed_3 <= RIN_M_CTRL_PC31DOWNTO12_intermed_2;
		RIN_M_CTRL_PC31DOWNTO12_intermed_4 <= RIN_M_CTRL_PC31DOWNTO12_intermed_3;
		RIN_M_CTRL_PC31DOWNTO12_intermed_5 <= RIN_M_CTRL_PC31DOWNTO12_intermed_4;
		IR_ADDR31DOWNTO12_intermed_1 <= IR.ADDR( 31 DOWNTO 12 );
		IR_ADDR31DOWNTO12_intermed_2 <= IR_ADDR31DOWNTO12_intermed_1;
		R_X_CTRL_PC31DOWNTO12_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 12 );
		R_X_CTRL_PC31DOWNTO12_intermed_2 <= R_X_CTRL_PC31DOWNTO12_intermed_1;
		R_X_CTRL_PC31DOWNTO12_intermed_3 <= R_X_CTRL_PC31DOWNTO12_intermed_2;
		V_D_PC31DOWNTO12_shadow_intermed_1 <= V_D_PC31DOWNTO12_shadow;
		V_D_PC31DOWNTO12_shadow_intermed_2 <= V_D_PC31DOWNTO12_shadow_intermed_1;
		V_D_PC31DOWNTO12_shadow_intermed_3 <= V_D_PC31DOWNTO12_shadow_intermed_2;
		V_D_PC31DOWNTO12_shadow_intermed_4 <= V_D_PC31DOWNTO12_shadow_intermed_3;
		V_D_PC31DOWNTO12_shadow_intermed_5 <= V_D_PC31DOWNTO12_shadow_intermed_4;
		V_D_PC31DOWNTO12_shadow_intermed_6 <= V_D_PC31DOWNTO12_shadow_intermed_5;
		V_D_PC31DOWNTO12_shadow_intermed_7 <= V_D_PC31DOWNTO12_shadow_intermed_6;
		V_D_PC31DOWNTO12_shadow_intermed_8 <= V_D_PC31DOWNTO12_shadow_intermed_7;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO12_shadow;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_4;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_6 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_5;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_7 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_6;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO12_shadow;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_3;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_5 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_4;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_6 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_5;
		EX_ADD_RES32DOWNTO330DOWNTO11_shadow_intermed_1 <= EX_ADD_RES32DOWNTO330DOWNTO11_shadow;
		EX_ADD_RES32DOWNTO330DOWNTO11_shadow_intermed_2 <= EX_ADD_RES32DOWNTO330DOWNTO11_shadow_intermed_1;
		RIN_F_PC31DOWNTO12_intermed_1 <= RIN.F.PC( 31 DOWNTO 12 );
		RIN_F_PC31DOWNTO12_intermed_2 <= RIN_F_PC31DOWNTO12_intermed_1;
		R_D_PC31DOWNTO12_intermed_1 <= R.D.PC( 31 DOWNTO 12 );
		R_D_PC31DOWNTO12_intermed_2 <= R_D_PC31DOWNTO12_intermed_1;
		R_D_PC31DOWNTO12_intermed_3 <= R_D_PC31DOWNTO12_intermed_2;
		R_D_PC31DOWNTO12_intermed_4 <= R_D_PC31DOWNTO12_intermed_3;
		R_D_PC31DOWNTO12_intermed_5 <= R_D_PC31DOWNTO12_intermed_4;
		R_D_PC31DOWNTO12_intermed_6 <= R_D_PC31DOWNTO12_intermed_5;
		R_D_PC31DOWNTO12_intermed_7 <= R_D_PC31DOWNTO12_intermed_6;
		R_A_CTRL_PC31DOWNTO12_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 12 );
		R_A_CTRL_PC31DOWNTO12_intermed_2 <= R_A_CTRL_PC31DOWNTO12_intermed_1;
		R_A_CTRL_PC31DOWNTO12_intermed_3 <= R_A_CTRL_PC31DOWNTO12_intermed_2;
		R_A_CTRL_PC31DOWNTO12_intermed_4 <= R_A_CTRL_PC31DOWNTO12_intermed_3;
		R_A_CTRL_PC31DOWNTO12_intermed_5 <= R_A_CTRL_PC31DOWNTO12_intermed_4;
		R_A_CTRL_PC31DOWNTO12_intermed_6 <= R_A_CTRL_PC31DOWNTO12_intermed_5;
		R_E_CTRL_PC31DOWNTO12_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 12 );
		R_E_CTRL_PC31DOWNTO12_intermed_2 <= R_E_CTRL_PC31DOWNTO12_intermed_1;
		R_E_CTRL_PC31DOWNTO12_intermed_3 <= R_E_CTRL_PC31DOWNTO12_intermed_2;
		R_E_CTRL_PC31DOWNTO12_intermed_4 <= R_E_CTRL_PC31DOWNTO12_intermed_3;
		R_E_CTRL_PC31DOWNTO12_intermed_5 <= R_E_CTRL_PC31DOWNTO12_intermed_4;
		RIN_X_CTRL_PC31DOWNTO12_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 12 );
		RIN_X_CTRL_PC31DOWNTO12_intermed_2 <= RIN_X_CTRL_PC31DOWNTO12_intermed_1;
		RIN_X_CTRL_PC31DOWNTO12_intermed_3 <= RIN_X_CTRL_PC31DOWNTO12_intermed_2;
		RIN_X_CTRL_PC31DOWNTO12_intermed_4 <= RIN_X_CTRL_PC31DOWNTO12_intermed_3;
		RIN_D_PC31DOWNTO12_intermed_1 <= RIN.D.PC( 31 DOWNTO 12 );
		RIN_D_PC31DOWNTO12_intermed_2 <= RIN_D_PC31DOWNTO12_intermed_1;
		RIN_D_PC31DOWNTO12_intermed_3 <= RIN_D_PC31DOWNTO12_intermed_2;
		RIN_D_PC31DOWNTO12_intermed_4 <= RIN_D_PC31DOWNTO12_intermed_3;
		RIN_D_PC31DOWNTO12_intermed_5 <= RIN_D_PC31DOWNTO12_intermed_4;
		RIN_D_PC31DOWNTO12_intermed_6 <= RIN_D_PC31DOWNTO12_intermed_5;
		RIN_D_PC31DOWNTO12_intermed_7 <= RIN_D_PC31DOWNTO12_intermed_6;
		RIN_D_PC31DOWNTO12_intermed_8 <= RIN_D_PC31DOWNTO12_intermed_7;
		VIR_ADDR31DOWNTO12_shadow_intermed_1 <= VIR_ADDR31DOWNTO12_shadow;
		VIR_ADDR31DOWNTO12_shadow_intermed_2 <= VIR_ADDR31DOWNTO12_shadow_intermed_1;
		VIR_ADDR31DOWNTO12_shadow_intermed_3 <= VIR_ADDR31DOWNTO12_shadow_intermed_2;
		V_F_PC31DOWNTO12_shadow_intermed_1 <= V_F_PC31DOWNTO12_shadow;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO12_shadow;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_4 <= V_M_CTRL_PC31DOWNTO12_shadow_intermed_3;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_5 <= V_M_CTRL_PC31DOWNTO12_shadow_intermed_4;
		ICO_DATA0_intermed_1 <= ICO.DATA ( 0 );
		RIN_D_INST0_intermed_1 <= RIN.D.INST ( 0 );
		V_D_INST0_shadow_intermed_1 <= V_D_INST0_shadow;
		V_D_INST0_shadow_intermed_2 <= V_D_INST0_shadow_intermed_1;
		R_D_INST0_intermed_1 <= R.D.INST( 0 );
		R_D_INST0_intermed_2 <= R_D_INST0_intermed_1;
		RIN_D_INST0_intermed_1 <= RIN.D.INST( 0 );
		RIN_D_INST0_intermed_2 <= RIN_D_INST0_intermed_1;
		V_D_INST0_shadow_intermed_1 <= V_D_INST0_shadow;
		V_D_INST1_shadow_intermed_1 <= V_D_INST1_shadow;
		V_D_INST1_shadow_intermed_2 <= V_D_INST1_shadow_intermed_1;
		RIN_D_INST1_intermed_1 <= RIN.D.INST ( 1 );
		RIN_D_INST1_intermed_1 <= RIN.D.INST( 1 );
		RIN_D_INST1_intermed_2 <= RIN_D_INST1_intermed_1;
		V_D_INST1_shadow_intermed_1 <= V_D_INST1_shadow;
		R_D_INST1_intermed_1 <= R.D.INST( 1 );
		R_D_INST1_intermed_2 <= R_D_INST1_intermed_1;
		ICO_DATA1_intermed_1 <= ICO.DATA ( 1 );
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA ( 0 )( 31 );
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_2 <= V_X_DATA031_shadow_intermed_1;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA( 0 )( 31 );
		RIN_X_DATA031_intermed_2 <= RIN_X_DATA031_intermed_1;
		DCO_DATA031_intermed_1 <= DCO.DATA ( 0 )( 31 );
		R_X_DATA031_intermed_1 <= R.X.DATA( 0 )( 31 );
		R_X_DATA031_intermed_2 <= R_X_DATA031_intermed_1;
		V_X_DATA1_shadow_intermed_1 <= V_X_DATA1_shadow;
		R_X_DATA1_intermed_1 <= R.X.DATA( 1 );
		RIN_X_DATA1_intermed_1 <= RIN.X.DATA( 1 );
		RIN_X_DATA1_intermed_2 <= RIN_X_DATA1_intermed_1;
		EX_JUMP_ADDRESS31DOWNTO12_shadow_intermed_1 <= EX_JUMP_ADDRESS31DOWNTO12_shadow;
		RIN_A_CTRL_PC31DOWNTO12_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 12 );
		RIN_A_CTRL_PC31DOWNTO12_intermed_2 <= RIN_A_CTRL_PC31DOWNTO12_intermed_1;
		RIN_A_CTRL_PC31DOWNTO12_intermed_3 <= RIN_A_CTRL_PC31DOWNTO12_intermed_2;
		RIN_A_CTRL_PC31DOWNTO12_intermed_4 <= RIN_A_CTRL_PC31DOWNTO12_intermed_3;
		RIN_A_CTRL_PC31DOWNTO12_intermed_5 <= RIN_A_CTRL_PC31DOWNTO12_intermed_4;
		RIN_A_CTRL_PC31DOWNTO12_intermed_6 <= RIN_A_CTRL_PC31DOWNTO12_intermed_5;
		RIN_E_CTRL_PC31DOWNTO12_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 12 );
		RIN_E_CTRL_PC31DOWNTO12_intermed_2 <= RIN_E_CTRL_PC31DOWNTO12_intermed_1;
		RIN_E_CTRL_PC31DOWNTO12_intermed_3 <= RIN_E_CTRL_PC31DOWNTO12_intermed_2;
		RIN_E_CTRL_PC31DOWNTO12_intermed_4 <= RIN_E_CTRL_PC31DOWNTO12_intermed_3;
		RIN_E_CTRL_PC31DOWNTO12_intermed_5 <= RIN_E_CTRL_PC31DOWNTO12_intermed_4;
		V_F_PC31DOWNTO12_shadow_intermed_1 <= V_F_PC31DOWNTO12_shadow;
		R_M_CTRL_PC31DOWNTO12_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 12 );
		R_M_CTRL_PC31DOWNTO12_intermed_2 <= R_M_CTRL_PC31DOWNTO12_intermed_1;
		R_M_CTRL_PC31DOWNTO12_intermed_3 <= R_M_CTRL_PC31DOWNTO12_intermed_2;
		IRIN_ADDR31DOWNTO12_intermed_1 <= IRIN.ADDR( 31 DOWNTO 12 );
		IRIN_ADDR31DOWNTO12_intermed_2 <= IRIN_ADDR31DOWNTO12_intermed_1;
		V_X_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO12_shadow;
		V_X_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_X_CTRL_PC31DOWNTO12_shadow_intermed_2;
		EX_ADD_RES32DOWNTO332DOWNTO13_shadow_intermed_1 <= EX_ADD_RES32DOWNTO332DOWNTO13_shadow;
		XC_TRAP_ADDRESS31DOWNTO12_shadow_intermed_1 <= XC_TRAP_ADDRESS31DOWNTO12_shadow;
		R_F_PC31DOWNTO12_intermed_1 <= R.F.PC( 31 DOWNTO 12 );
		RIN_M_CTRL_PC31DOWNTO12_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 12 );
		RIN_M_CTRL_PC31DOWNTO12_intermed_2 <= RIN_M_CTRL_PC31DOWNTO12_intermed_1;
		RIN_M_CTRL_PC31DOWNTO12_intermed_3 <= RIN_M_CTRL_PC31DOWNTO12_intermed_2;
		RIN_M_CTRL_PC31DOWNTO12_intermed_4 <= RIN_M_CTRL_PC31DOWNTO12_intermed_3;
		IR_ADDR31DOWNTO12_intermed_1 <= IR.ADDR( 31 DOWNTO 12 );
		R_X_CTRL_PC31DOWNTO12_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 12 );
		R_X_CTRL_PC31DOWNTO12_intermed_2 <= R_X_CTRL_PC31DOWNTO12_intermed_1;
		V_D_PC31DOWNTO12_shadow_intermed_1 <= V_D_PC31DOWNTO12_shadow;
		V_D_PC31DOWNTO12_shadow_intermed_2 <= V_D_PC31DOWNTO12_shadow_intermed_1;
		V_D_PC31DOWNTO12_shadow_intermed_3 <= V_D_PC31DOWNTO12_shadow_intermed_2;
		V_D_PC31DOWNTO12_shadow_intermed_4 <= V_D_PC31DOWNTO12_shadow_intermed_3;
		V_D_PC31DOWNTO12_shadow_intermed_5 <= V_D_PC31DOWNTO12_shadow_intermed_4;
		V_D_PC31DOWNTO12_shadow_intermed_6 <= V_D_PC31DOWNTO12_shadow_intermed_5;
		V_D_PC31DOWNTO12_shadow_intermed_7 <= V_D_PC31DOWNTO12_shadow_intermed_6;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO12_shadow;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_4;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_6 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_5;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO12_shadow;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_3;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_5 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_4;
		EX_ADD_RES32DOWNTO330DOWNTO11_shadow_intermed_1 <= EX_ADD_RES32DOWNTO330DOWNTO11_shadow;
		RIN_F_PC31DOWNTO12_intermed_1 <= RIN.F.PC( 31 DOWNTO 12 );
		RIN_F_PC31DOWNTO12_intermed_2 <= RIN_F_PC31DOWNTO12_intermed_1;
		R_D_PC31DOWNTO12_intermed_1 <= R.D.PC( 31 DOWNTO 12 );
		R_D_PC31DOWNTO12_intermed_2 <= R_D_PC31DOWNTO12_intermed_1;
		R_D_PC31DOWNTO12_intermed_3 <= R_D_PC31DOWNTO12_intermed_2;
		R_D_PC31DOWNTO12_intermed_4 <= R_D_PC31DOWNTO12_intermed_3;
		R_D_PC31DOWNTO12_intermed_5 <= R_D_PC31DOWNTO12_intermed_4;
		R_D_PC31DOWNTO12_intermed_6 <= R_D_PC31DOWNTO12_intermed_5;
		R_A_CTRL_PC31DOWNTO12_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 12 );
		R_A_CTRL_PC31DOWNTO12_intermed_2 <= R_A_CTRL_PC31DOWNTO12_intermed_1;
		R_A_CTRL_PC31DOWNTO12_intermed_3 <= R_A_CTRL_PC31DOWNTO12_intermed_2;
		R_A_CTRL_PC31DOWNTO12_intermed_4 <= R_A_CTRL_PC31DOWNTO12_intermed_3;
		R_A_CTRL_PC31DOWNTO12_intermed_5 <= R_A_CTRL_PC31DOWNTO12_intermed_4;
		R_E_CTRL_PC31DOWNTO12_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 12 );
		R_E_CTRL_PC31DOWNTO12_intermed_2 <= R_E_CTRL_PC31DOWNTO12_intermed_1;
		R_E_CTRL_PC31DOWNTO12_intermed_3 <= R_E_CTRL_PC31DOWNTO12_intermed_2;
		R_E_CTRL_PC31DOWNTO12_intermed_4 <= R_E_CTRL_PC31DOWNTO12_intermed_3;
		RIN_X_CTRL_PC31DOWNTO12_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 12 );
		RIN_X_CTRL_PC31DOWNTO12_intermed_2 <= RIN_X_CTRL_PC31DOWNTO12_intermed_1;
		RIN_X_CTRL_PC31DOWNTO12_intermed_3 <= RIN_X_CTRL_PC31DOWNTO12_intermed_2;
		RIN_D_PC31DOWNTO12_intermed_1 <= RIN.D.PC( 31 DOWNTO 12 );
		RIN_D_PC31DOWNTO12_intermed_2 <= RIN_D_PC31DOWNTO12_intermed_1;
		RIN_D_PC31DOWNTO12_intermed_3 <= RIN_D_PC31DOWNTO12_intermed_2;
		RIN_D_PC31DOWNTO12_intermed_4 <= RIN_D_PC31DOWNTO12_intermed_3;
		RIN_D_PC31DOWNTO12_intermed_5 <= RIN_D_PC31DOWNTO12_intermed_4;
		RIN_D_PC31DOWNTO12_intermed_6 <= RIN_D_PC31DOWNTO12_intermed_5;
		RIN_D_PC31DOWNTO12_intermed_7 <= RIN_D_PC31DOWNTO12_intermed_6;
		VIR_ADDR31DOWNTO12_shadow_intermed_1 <= VIR_ADDR31DOWNTO12_shadow;
		VIR_ADDR31DOWNTO12_shadow_intermed_2 <= VIR_ADDR31DOWNTO12_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO12_shadow;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_4 <= V_M_CTRL_PC31DOWNTO12_shadow_intermed_3;
		V_D_INST0_shadow_intermed_1 <= V_D_INST0_shadow;
		R_D_INST0_intermed_1 <= R.D.INST( 0 );
		RIN_D_INST0_intermed_1 <= RIN.D.INST( 0 );
		RIN_D_INST0_intermed_2 <= RIN_D_INST0_intermed_1;
		V_D_INST1_shadow_intermed_1 <= V_D_INST1_shadow;
		RIN_D_INST1_intermed_1 <= RIN.D.INST( 1 );
		RIN_D_INST1_intermed_2 <= RIN_D_INST1_intermed_1;
		R_D_INST1_intermed_1 <= R.D.INST( 1 );
		V_X_DATA03_shadow_intermed_1 <= V_X_DATA03_shadow;
		V_X_DATA03_shadow_intermed_2 <= V_X_DATA03_shadow_intermed_1;
		V_X_DATA03_shadow_intermed_1 <= V_X_DATA03_shadow;
		DCO_DATA03_intermed_1 <= DCO.DATA ( 0 )( 3 );
		RIN_X_DATA03_intermed_1 <= RIN.X.DATA ( 0 )( 3 );
		R_X_DATA03_intermed_1 <= R.X.DATA( 0 )( 3 );
		R_X_DATA03_intermed_2 <= R_X_DATA03_intermed_1;
		RIN_X_DATA03_intermed_1 <= RIN.X.DATA( 0 )( 3 );
		RIN_X_DATA03_intermed_2 <= RIN_X_DATA03_intermed_1;
		V_X_DATA03_shadow_intermed_1 <= V_X_DATA03_shadow;
		R_X_DATA03_intermed_1 <= R.X.DATA( 0 )( 3 );
		RIN_X_DATA03_intermed_1 <= RIN.X.DATA( 0 )( 3 );
		RIN_X_DATA03_intermed_2 <= RIN_X_DATA03_intermed_1;
		V_A_CTRL_INST20_shadow_intermed_1 <= V_A_CTRL_INST20_shadow;
		RIN_A_CTRL_INST20_intermed_1 <= RIN.A.CTRL.INST ( 20 );
		RIN_A_CTRL_INST20_intermed_1 <= RIN.A.CTRL.INST( 20 );
		RIN_A_CTRL_INST20_intermed_2 <= RIN_A_CTRL_INST20_intermed_1;
		DE_INST20_shadow_intermed_1 <= DE_INST20_shadow;
		DE_INST20_shadow_intermed_2 <= DE_INST20_shadow_intermed_1;
		V_A_CTRL_INST20_shadow_intermed_1 <= V_A_CTRL_INST20_shadow;
		V_A_CTRL_INST20_shadow_intermed_2 <= V_A_CTRL_INST20_shadow_intermed_1;
		R_A_CTRL_INST20_intermed_1 <= R.A.CTRL.INST( 20 );
		R_A_CTRL_INST20_intermed_2 <= R_A_CTRL_INST20_intermed_1;
		RIN_X_DATA00_intermed_1 <= RIN.X.DATA ( 0 )( 0 );
		DCO_DATA00_intermed_1 <= DCO.DATA ( 0 )( 0 );
		V_X_DATA00_shadow_intermed_1 <= V_X_DATA00_shadow;
		V_X_DATA00_shadow_intermed_1 <= V_X_DATA00_shadow;
		V_X_DATA00_shadow_intermed_2 <= V_X_DATA00_shadow_intermed_1;
		RIN_X_DATA00_intermed_1 <= RIN.X.DATA( 0 )( 0 );
		RIN_X_DATA00_intermed_2 <= RIN_X_DATA00_intermed_1;
		R_X_DATA00_intermed_1 <= R.X.DATA( 0 )( 0 );
		R_X_DATA00_intermed_2 <= R_X_DATA00_intermed_1;
		V_X_DATA04DOWNTO0_shadow_intermed_1 <= V_X_DATA04DOWNTO0_shadow;
		V_X_DATA04DOWNTO0_shadow_intermed_2 <= V_X_DATA04DOWNTO0_shadow_intermed_1;
		R_X_DATA04DOWNTO0_intermed_1 <= R.X.DATA( 0 )( 4 DOWNTO 0 );
		R_X_DATA04DOWNTO0_intermed_2 <= R_X_DATA04DOWNTO0_intermed_1;
		DCO_DATA04DOWNTO0_intermed_1 <= DCO.DATA ( 0 )( 4 DOWNTO 0 );
		RIN_X_DATA04DOWNTO0_intermed_1 <= RIN.X.DATA( 0 )( 4 DOWNTO 0 );
		RIN_X_DATA04DOWNTO0_intermed_2 <= RIN_X_DATA04DOWNTO0_intermed_1;
		RIN_X_DATA04DOWNTO0_intermed_1 <= RIN.X.DATA ( 0 )( 4 DOWNTO 0 );
		V_X_DATA04DOWNTO0_shadow_intermed_1 <= V_X_DATA04DOWNTO0_shadow;
		V_A_CTRL_INST24_shadow_intermed_1 <= V_A_CTRL_INST24_shadow;
		V_A_CTRL_INST24_shadow_intermed_2 <= V_A_CTRL_INST24_shadow_intermed_1;
		DE_INST24_shadow_intermed_1 <= DE_INST24_shadow;
		DE_INST24_shadow_intermed_2 <= DE_INST24_shadow_intermed_1;
		R_A_CTRL_INST24_intermed_1 <= R.A.CTRL.INST( 24 );
		R_A_CTRL_INST24_intermed_2 <= R_A_CTRL_INST24_intermed_1;
		RIN_A_CTRL_INST24_intermed_1 <= RIN.A.CTRL.INST ( 24 );
		V_A_CTRL_INST24_shadow_intermed_1 <= V_A_CTRL_INST24_shadow;
		RIN_A_CTRL_INST24_intermed_1 <= RIN.A.CTRL.INST( 24 );
		RIN_A_CTRL_INST24_intermed_2 <= RIN_A_CTRL_INST24_intermed_1;
		RIN_A_CTRL_INST20_intermed_1 <= RIN.A.CTRL.INST( 20 );
		RIN_A_CTRL_INST20_intermed_2 <= RIN_A_CTRL_INST20_intermed_1;
		DE_INST20_shadow_intermed_1 <= DE_INST20_shadow;
		V_A_CTRL_INST20_shadow_intermed_1 <= V_A_CTRL_INST20_shadow;
		R_A_CTRL_INST20_intermed_1 <= R.A.CTRL.INST( 20 );
		V_A_CTRL_INST24_shadow_intermed_1 <= V_A_CTRL_INST24_shadow;
		DE_INST24_shadow_intermed_1 <= DE_INST24_shadow;
		R_A_CTRL_INST24_intermed_1 <= R.A.CTRL.INST( 24 );
		RIN_A_CTRL_INST24_intermed_1 <= RIN.A.CTRL.INST( 24 );
		RIN_A_CTRL_INST24_intermed_2 <= RIN_A_CTRL_INST24_intermed_1;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1;
		R_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= R.X.RESULT( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		R_X_RESULT6DOWNTO03DOWNTO0_intermed_2 <= R_X_RESULT6DOWNTO03DOWNTO0_intermed_1;
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= RIN.X.RESULT( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2 <= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1;
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= RIN.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow;
		R_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= R.X.RESULT( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= RIN.X.RESULT( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2 <= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1;
		RIN_F_PC_intermed_1 <= RIN.F.PC;
		EX_ADD_RES32DOWNTO3_shadow_intermed_1 <= EX_ADD_RES32DOWNTO3_shadow;
		XC_TRAP_ADDRESS_shadow_intermed_1 <= XC_TRAP_ADDRESS_shadow;
		EX_JUMP_ADDRESS_shadow_intermed_1 <= EX_JUMP_ADDRESS_shadow;
		V_F_PC_shadow_intermed_1 <= V_F_PC_shadow;
		RIN_A_RFE1_intermed_1 <= RIN.A.RFE1;
		V_A_RFE1_shadow_intermed_1 <= V_A_RFE1_shadow;
		RIN_A_RFE2_intermed_1 <= RIN.A.RFE2;
		V_A_RFE2_shadow_intermed_1 <= V_A_RFE2_shadow;
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		V_X_DATA0_shadow_intermed_2 <= V_X_DATA0_shadow_intermed_1;
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA ( 0 );
		V_E_OP1_shadow_intermed_1 <= V_E_OP1_shadow;
		V_E_OP2_shadow_intermed_1 <= V_E_OP2_shadow;
		RIN_E_OP2_intermed_1 <= RIN.E.OP2;
		RIN_E_OP1_intermed_1 <= RIN.E.OP1;
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		V_E_ALUCIN_shadow_intermed_1 <= V_E_ALUCIN_shadow;
		R_X_DATA0_intermed_1 <= R.X.DATA( 0 );
		RIN_E_ALUCIN_intermed_1 <= RIN.E.ALUCIN;
		DCO_DATA0_intermed_1 <= DCO.DATA ( 0 );
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA( 0 );
		RIN_X_DATA0_intermed_2 <= RIN_X_DATA0_intermed_1;
		RIN_X_DATA00_intermed_1 <= RIN.X.DATA ( 0 )( 0 );
		RIN_X_DATA00_intermed_2 <= RIN_X_DATA00_intermed_1;
		V_X_DATA00_shadow_intermed_1 <= V_X_DATA00_shadow;
		DCO_DATA00_intermed_1 <= DCO.DATA ( 0 )( 0 );
		V_X_DATA00_shadow_intermed_1 <= V_X_DATA00_shadow;
		V_X_DATA00_shadow_intermed_2 <= V_X_DATA00_shadow_intermed_1;
		V_E_YMSB_shadow_intermed_1 <= V_E_YMSB_shadow;
		RIN_X_DATA00_intermed_1 <= RIN.X.DATA ( 0 ) ( 0 );
		V_X_DATA00_shadow_intermed_1 <= V_X_DATA00_shadow;
		V_X_DATA00_shadow_intermed_2 <= V_X_DATA00_shadow_intermed_1;
		V_X_DATA00_shadow_intermed_3 <= V_X_DATA00_shadow_intermed_2;
		R_X_DATA00_intermed_1 <= R.X.DATA ( 0 )( 0 );
		RIN_X_DATA00_intermed_1 <= RIN.X.DATA( 0 )( 0 );
		RIN_X_DATA00_intermed_2 <= RIN_X_DATA00_intermed_1;
		RIN_X_DATA00_intermed_3 <= RIN_X_DATA00_intermed_2;
		R_X_DATA00_intermed_1 <= R.X.DATA( 0 )( 0 );
		R_X_DATA00_intermed_2 <= R_X_DATA00_intermed_1;
		RIN_E_YMSB_intermed_1 <= RIN.E.YMSB;
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		V_X_DATA0_shadow_intermed_2 <= V_X_DATA0_shadow_intermed_1;
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA ( 0 );
		V_E_OP1_shadow_intermed_1 <= V_E_OP1_shadow;
		RIN_E_OP1_intermed_1 <= RIN.E.OP1;
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		R_X_DATA0_intermed_1 <= R.X.DATA( 0 );
		DCO_DATA0_intermed_1 <= DCO.DATA ( 0 );
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA( 0 );
		RIN_X_DATA0_intermed_2 <= RIN_X_DATA0_intermed_1;
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		V_X_DATA0_shadow_intermed_2 <= V_X_DATA0_shadow_intermed_1;
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA ( 0 );
		V_E_OP2_shadow_intermed_1 <= V_E_OP2_shadow;
		RIN_E_OP2_intermed_1 <= RIN.E.OP2;
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		R_X_DATA0_intermed_1 <= R.X.DATA( 0 );
		DCO_DATA0_intermed_1 <= DCO.DATA ( 0 );
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA( 0 );
		RIN_X_DATA0_intermed_2 <= RIN_X_DATA0_intermed_1;
		RIN_X_DATA04DOWNTO0_intermed_1 <= RIN.X.DATA ( 0 ) ( 4 DOWNTO 0 );
		V_X_DATA04DOWNTO0_shadow_intermed_1 <= V_X_DATA04DOWNTO0_shadow;
		V_X_DATA04DOWNTO0_shadow_intermed_2 <= V_X_DATA04DOWNTO0_shadow_intermed_1;
		V_X_DATA04DOWNTO0_shadow_intermed_3 <= V_X_DATA04DOWNTO0_shadow_intermed_2;
		R_X_DATA04DOWNTO0_intermed_1 <= R.X.DATA( 0 )( 4 DOWNTO 0 );
		R_X_DATA04DOWNTO0_intermed_2 <= R_X_DATA04DOWNTO0_intermed_1;
		V_E_SHCNT_shadow_intermed_1 <= V_E_SHCNT_shadow;
		R_X_DATA04DOWNTO0_intermed_1 <= R.X.DATA ( 0 )( 4 DOWNTO 0 );
		V_X_DATA04DOWNTO0_shadow_intermed_1 <= V_X_DATA04DOWNTO0_shadow;
		RIN_X_DATA04DOWNTO0_intermed_1 <= RIN.X.DATA( 0 )( 4 DOWNTO 0 );
		RIN_X_DATA04DOWNTO0_intermed_2 <= RIN_X_DATA04DOWNTO0_intermed_1;
		RIN_X_DATA04DOWNTO0_intermed_3 <= RIN_X_DATA04DOWNTO0_intermed_2;
		RIN_X_DATA04DOWNTO0_intermed_1 <= RIN.X.DATA ( 0 )( 4 DOWNTO 0 );
		RIN_X_DATA04DOWNTO0_intermed_2 <= RIN_X_DATA04DOWNTO0_intermed_1;
		DCO_DATA04DOWNTO0_intermed_1 <= DCO.DATA ( 0 )( 4 DOWNTO 0 );
		RIN_E_SHCNT_intermed_1 <= RIN.E.SHCNT;
		V_X_DATA04DOWNTO0_shadow_intermed_1 <= V_X_DATA04DOWNTO0_shadow;
		V_X_DATA04DOWNTO0_shadow_intermed_2 <= V_X_DATA04DOWNTO0_shadow_intermed_1;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA ( 0 )( 31 );
		RIN_X_DATA031_intermed_2 <= RIN_X_DATA031_intermed_1;
		DE_INST19_shadow_intermed_1 <= DE_INST19_shadow;
		DE_INST19_shadow_intermed_2 <= DE_INST19_shadow_intermed_1;
		V_A_CTRL_INST20_shadow_intermed_1 <= V_A_CTRL_INST20_shadow;
		V_A_CTRL_INST20_shadow_intermed_2 <= V_A_CTRL_INST20_shadow_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_3 <= V_A_CTRL_INST19_shadow_intermed_2;
		RIN_A_CTRL_INST20_intermed_1 <= RIN.A.CTRL.INST ( 20 );
		RIN_A_CTRL_INST20_intermed_2 <= RIN_A_CTRL_INST20_intermed_1;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_2 <= V_X_DATA031_shadow_intermed_1;
		V_E_CTRL_INST19_shadow_intermed_1 <= V_E_CTRL_INST19_shadow;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_2 <= V_X_DATA031_shadow_intermed_1;
		V_X_DATA031_shadow_intermed_3 <= V_X_DATA031_shadow_intermed_2;
		V_E_CTRL_INST19_shadow_intermed_1 <= V_E_CTRL_INST19_shadow;
		V_E_CTRL_INST19_shadow_intermed_2 <= V_E_CTRL_INST19_shadow_intermed_1;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA( 0 )( 31 );
		RIN_X_DATA031_intermed_2 <= RIN_X_DATA031_intermed_1;
		RIN_X_DATA031_intermed_3 <= RIN_X_DATA031_intermed_2;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA ( 0 ) ( 31 );
		V_E_SARI_shadow_intermed_1 <= V_E_SARI_shadow;
		R_E_CTRL_INST19_intermed_1 <= R.E.CTRL.INST( 19 );
		DCO_DATA031_intermed_1 <= DCO.DATA ( 0 )( 31 );
		R_X_DATA031_intermed_1 <= R.X.DATA( 0 )( 31 );
		R_X_DATA031_intermed_2 <= R_X_DATA031_intermed_1;
		RIN_E_CTRL_INST20_intermed_1 <= RIN.E.CTRL.INST ( 20 );
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST ( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		R_E_CTRL_INST20_intermed_1 <= R.E.CTRL.INST( 20 );
		R_A_CTRL_INST20_intermed_1 <= R.A.CTRL.INST ( 20 );
		RIN_A_CTRL_INST20_intermed_1 <= RIN.A.CTRL.INST( 20 );
		RIN_A_CTRL_INST20_intermed_2 <= RIN_A_CTRL_INST20_intermed_1;
		RIN_A_CTRL_INST20_intermed_3 <= RIN_A_CTRL_INST20_intermed_2;
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST( 19 );
		R_A_CTRL_INST19_intermed_2 <= R_A_CTRL_INST19_intermed_1;
		V_E_CTRL_INST20_shadow_intermed_1 <= V_E_CTRL_INST20_shadow;
		V_E_CTRL_INST20_shadow_intermed_2 <= V_E_CTRL_INST20_shadow_intermed_1;
		V_E_CTRL_INST20_shadow_intermed_1 <= V_E_CTRL_INST20_shadow;
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST ( 19 );
		DE_INST20_shadow_intermed_1 <= DE_INST20_shadow;
		DE_INST20_shadow_intermed_2 <= DE_INST20_shadow_intermed_1;
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		RIN_A_CTRL_INST19_intermed_3 <= RIN_A_CTRL_INST19_intermed_2;
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST ( 19 );
		V_A_CTRL_INST20_shadow_intermed_1 <= V_A_CTRL_INST20_shadow;
		V_A_CTRL_INST20_shadow_intermed_2 <= V_A_CTRL_INST20_shadow_intermed_1;
		V_A_CTRL_INST20_shadow_intermed_3 <= V_A_CTRL_INST20_shadow_intermed_2;
		R_X_DATA031_intermed_1 <= R.X.DATA ( 0 )( 31 );
		RIN_E_SARI_intermed_1 <= RIN.E.SARI;
		RIN_E_CTRL_INST20_intermed_1 <= RIN.E.CTRL.INST( 20 );
		RIN_E_CTRL_INST20_intermed_2 <= RIN_E_CTRL_INST20_intermed_1;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST( 19 );
		RIN_E_CTRL_INST19_intermed_2 <= RIN_E_CTRL_INST19_intermed_1;
		R_A_CTRL_INST20_intermed_1 <= R.A.CTRL.INST( 20 );
		R_A_CTRL_INST20_intermed_2 <= R_A_CTRL_INST20_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		V_M_DCI_SIGNED_shadow_intermed_1 <= V_M_DCI_SIGNED_shadow;
		V_M_DCI_SIGNED_shadow_intermed_2 <= V_M_DCI_SIGNED_shadow_intermed_1;
		RIN_M_DCI_SIGNED_intermed_1 <= RIN.M.DCI.SIGNED;
		RIN_M_DCI_SIGNED_intermed_2 <= RIN_M_DCI_SIGNED_intermed_1;
		R_M_DCI_SIGNED_intermed_1 <= R.M.DCI.SIGNED;
		V_X_DCI_SIGNED_shadow_intermed_1 <= V_X_DCI_SIGNED_shadow;
		RIN_X_DCI_SIGNED_intermed_1 <= RIN.X.DCI.SIGNED;
		RIN_M_DCI_SIZE_intermed_1 <= RIN.M.DCI.SIZE;
		RIN_M_DCI_SIZE_intermed_2 <= RIN_M_DCI_SIZE_intermed_1;
		V_M_DCI_SIZE_shadow_intermed_1 <= V_M_DCI_SIZE_shadow;
		V_M_DCI_SIZE_shadow_intermed_2 <= V_M_DCI_SIZE_shadow_intermed_1;
		R_M_DCI_SIZE_intermed_1 <= R.M.DCI.SIZE;
		V_X_DCI_SIZE_shadow_intermed_1 <= V_X_DCI_SIZE_shadow;
		RIN_X_DCI_SIZE_intermed_1 <= RIN.X.DCI.SIZE;
		V_M_RESULT1DOWNTO0_shadow_intermed_1 <= V_M_RESULT1DOWNTO0_shadow;
		V_M_RESULT1DOWNTO0_shadow_intermed_2 <= V_M_RESULT1DOWNTO0_shadow_intermed_1;
		V_M_RESULT1DOWNTO0_shadow_intermed_3 <= V_M_RESULT1DOWNTO0_shadow_intermed_2;
		RIN_X_LADDR_intermed_1 <= RIN.X.LADDR;
		R_M_RESULT1DOWNTO0_intermed_1 <= R.M.RESULT ( 1 DOWNTO 0 );
		RIN_M_RESULT1DOWNTO0_intermed_1 <= RIN.M.RESULT ( 1 DOWNTO 0 );
		RIN_M_RESULT1DOWNTO0_intermed_2 <= RIN_M_RESULT1DOWNTO0_intermed_1;
		RIN_M_RESULT1DOWNTO0_intermed_1 <= RIN.M.RESULT( 1 DOWNTO 0 );
		RIN_M_RESULT1DOWNTO0_intermed_2 <= RIN_M_RESULT1DOWNTO0_intermed_1;
		RIN_M_RESULT1DOWNTO0_intermed_3 <= RIN_M_RESULT1DOWNTO0_intermed_2;
		V_M_RESULT1DOWNTO0_shadow_intermed_1 <= V_M_RESULT1DOWNTO0_shadow;
		V_M_RESULT1DOWNTO0_shadow_intermed_2 <= V_M_RESULT1DOWNTO0_shadow_intermed_1;
		V_X_LADDR_shadow_intermed_1 <= V_X_LADDR_shadow;
		R_M_RESULT1DOWNTO0_intermed_1 <= R.M.RESULT( 1 DOWNTO 0 );
		R_M_RESULT1DOWNTO0_intermed_2 <= R_M_RESULT1DOWNTO0_intermed_1;
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		V_X_DATA0_shadow_intermed_2 <= V_X_DATA0_shadow_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 2 );
		R_M_CTRL_PC31DOWNTO2_intermed_2 <= R_M_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_3 <= RIN_M_CTRL_PC31DOWNTO2_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		RIN_A_CTRL_PC31DOWNTO2_intermed_5 <= RIN_A_CTRL_PC31DOWNTO2_intermed_4;
		RIN_X_RESULT_intermed_1 <= RIN.X.RESULT;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO2_shadow;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_4 <= R_A_CTRL_PC31DOWNTO2_intermed_3;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2;
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA ( 0 );
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC ( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		V_X_RESULT_shadow_intermed_1 <= V_X_RESULT_shadow;
		R_X_CTRL_PC31DOWNTO2_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC ( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_5 <= V_D_PC31DOWNTO2_shadow_intermed_4;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_5 <= RIN_D_PC31DOWNTO2_intermed_4;
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC ( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC ( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC ( 31 DOWNTO 2 );
		R_X_DATA0_intermed_1 <= R.X.DATA( 0 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_2 <= RIN_X_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC ( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_3 <= R_E_CTRL_PC31DOWNTO2_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		R_D_PC31DOWNTO2_intermed_4 <= R_D_PC31DOWNTO2_intermed_3;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC ( 31 DOWNTO 2 );
		DCO_DATA0_intermed_1 <= DCO.DATA ( 0 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_4 <= RIN_E_CTRL_PC31DOWNTO2_intermed_3;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO2_shadow;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA( 0 );
		RIN_X_DATA0_intermed_2 <= RIN_X_DATA0_intermed_1;
		V_X_ANNUL_ALL_shadow_intermed_1 <= V_X_ANNUL_ALL_shadow;
		V_X_ANNUL_ALL_shadow_intermed_2 <= V_X_ANNUL_ALL_shadow_intermed_1;
		V_X_ANNUL_ALL_shadow_intermed_3 <= V_X_ANNUL_ALL_shadow_intermed_2;
		V_X_ANNUL_ALL_shadow_intermed_4 <= V_X_ANNUL_ALL_shadow_intermed_3;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_A_CTRL_ANNUL_intermed_2 <= RIN_A_CTRL_ANNUL_intermed_1;
		RIN_A_CTRL_ANNUL_intermed_3 <= RIN_A_CTRL_ANNUL_intermed_2;
		RIN_A_CTRL_ANNUL_intermed_4 <= RIN_A_CTRL_ANNUL_intermed_3;
		RIN_A_CTRL_ANNUL_intermed_5 <= RIN_A_CTRL_ANNUL_intermed_4;
		R_M_CTRL_WREG_intermed_1 <= R.M.CTRL.WREG;
		R_A_CTRL_ANNUL_intermed_1 <= R.A.CTRL.ANNUL;
		R_A_CTRL_ANNUL_intermed_2 <= R_A_CTRL_ANNUL_intermed_1;
		R_A_CTRL_ANNUL_intermed_3 <= R_A_CTRL_ANNUL_intermed_2;
		R_A_CTRL_ANNUL_intermed_4 <= R_A_CTRL_ANNUL_intermed_3;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_X_ANNUL_ALL_intermed_2 <= RIN_X_ANNUL_ALL_intermed_1;
		RIN_X_ANNUL_ALL_intermed_3 <= RIN_X_ANNUL_ALL_intermed_2;
		RIN_X_ANNUL_ALL_intermed_4 <= RIN_X_ANNUL_ALL_intermed_3;
		RIN_X_ANNUL_ALL_intermed_5 <= RIN_X_ANNUL_ALL_intermed_4;
		V_M_CTRL_WREG_shadow_intermed_1 <= V_M_CTRL_WREG_shadow;
		V_M_CTRL_WREG_shadow_intermed_2 <= V_M_CTRL_WREG_shadow_intermed_1;
		R_X_ANNUL_ALL_intermed_1 <= R.X.ANNUL_ALL;
		R_X_ANNUL_ALL_intermed_2 <= R_X_ANNUL_ALL_intermed_1;
		R_X_ANNUL_ALL_intermed_3 <= R_X_ANNUL_ALL_intermed_2;
		R_X_ANNUL_ALL_intermed_4 <= R_X_ANNUL_ALL_intermed_3;
		V_X_CTRL_WREG_shadow_intermed_1 <= V_X_CTRL_WREG_shadow;
		R_E_CTRL_WREG_intermed_1 <= R.E.CTRL.WREG;
		R_E_CTRL_WREG_intermed_2 <= R_E_CTRL_WREG_intermed_1;
		RIN_X_CTRL_WREG_intermed_1 <= RIN.X.CTRL.WREG;
		V_A_CTRL_ANNUL_shadow_intermed_1 <= V_A_CTRL_ANNUL_shadow;
		V_A_CTRL_ANNUL_shadow_intermed_2 <= V_A_CTRL_ANNUL_shadow_intermed_1;
		V_A_CTRL_ANNUL_shadow_intermed_3 <= V_A_CTRL_ANNUL_shadow_intermed_2;
		V_A_CTRL_ANNUL_shadow_intermed_4 <= V_A_CTRL_ANNUL_shadow_intermed_3;
		RIN_E_CTRL_WREG_intermed_1 <= RIN.E.CTRL.WREG;
		RIN_E_CTRL_WREG_intermed_2 <= RIN_E_CTRL_WREG_intermed_1;
		RIN_E_CTRL_WREG_intermed_3 <= RIN_E_CTRL_WREG_intermed_2;
		RIN_M_CTRL_WREG_intermed_1 <= RIN.M.CTRL.WREG;
		RIN_M_CTRL_WREG_intermed_2 <= RIN_M_CTRL_WREG_intermed_1;
		V_E_CTRL_WREG_shadow_intermed_1 <= V_E_CTRL_WREG_shadow;
		V_E_CTRL_WREG_shadow_intermed_2 <= V_E_CTRL_WREG_shadow_intermed_1;
		V_E_CTRL_WREG_shadow_intermed_3 <= V_E_CTRL_WREG_shadow_intermed_2;
		RIN_A_CTRL_WREG_intermed_1 <= RIN.A.CTRL.WREG;
		RIN_A_CTRL_WREG_intermed_2 <= RIN_A_CTRL_WREG_intermed_1;
		RIN_A_CTRL_WREG_intermed_3 <= RIN_A_CTRL_WREG_intermed_2;
		RIN_A_CTRL_WREG_intermed_4 <= RIN_A_CTRL_WREG_intermed_3;
		V_A_CTRL_WREG_shadow_intermed_1 <= V_A_CTRL_WREG_shadow;
		V_A_CTRL_WREG_shadow_intermed_2 <= V_A_CTRL_WREG_shadow_intermed_1;
		V_A_CTRL_WREG_shadow_intermed_3 <= V_A_CTRL_WREG_shadow_intermed_2;
		V_A_CTRL_WREG_shadow_intermed_4 <= V_A_CTRL_WREG_shadow_intermed_3;
		R_A_CTRL_WREG_intermed_1 <= R.A.CTRL.WREG;
		R_A_CTRL_WREG_intermed_2 <= R_A_CTRL_WREG_intermed_1;
		R_A_CTRL_WREG_intermed_3 <= R_A_CTRL_WREG_intermed_2;
		V_E_CTRL_TT_shadow_intermed_1 <= V_E_CTRL_TT_shadow;
		V_E_CTRL_TT_shadow_intermed_2 <= V_E_CTRL_TT_shadow_intermed_1;
		V_E_CTRL_TT_shadow_intermed_3 <= V_E_CTRL_TT_shadow_intermed_2;
		V_X_CTRL_TT_shadow_intermed_1 <= V_X_CTRL_TT_shadow;
		V_X_RESULT6DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO0_shadow;
		V_X_RESULT6DOWNTO0_shadow_intermed_2 <= V_X_RESULT6DOWNTO0_shadow_intermed_1;
		RIN_A_CTRL_TT_intermed_1 <= RIN.A.CTRL.TT;
		RIN_A_CTRL_TT_intermed_2 <= RIN_A_CTRL_TT_intermed_1;
		RIN_A_CTRL_TT_intermed_3 <= RIN_A_CTRL_TT_intermed_2;
		RIN_A_CTRL_TT_intermed_4 <= RIN_A_CTRL_TT_intermed_3;
		RIN_X_RESULT6DOWNTO0_intermed_1 <= RIN.X.RESULT( 6 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO0_intermed_2 <= RIN_X_RESULT6DOWNTO0_intermed_1;
		RIN_E_CTRL_TT_intermed_1 <= RIN.E.CTRL.TT;
		RIN_E_CTRL_TT_intermed_2 <= RIN_E_CTRL_TT_intermed_1;
		RIN_E_CTRL_TT_intermed_3 <= RIN_E_CTRL_TT_intermed_2;
		V_M_CTRL_TT_shadow_intermed_1 <= V_M_CTRL_TT_shadow;
		V_M_CTRL_TT_shadow_intermed_2 <= V_M_CTRL_TT_shadow_intermed_1;
		R_X_RESULT6DOWNTO0_intermed_1 <= R.X.RESULT( 6 DOWNTO 0 );
		R_A_CTRL_TT_intermed_1 <= R.A.CTRL.TT;
		R_A_CTRL_TT_intermed_2 <= R_A_CTRL_TT_intermed_1;
		R_A_CTRL_TT_intermed_3 <= R_A_CTRL_TT_intermed_2;
		V_A_CTRL_TT_shadow_intermed_1 <= V_A_CTRL_TT_shadow;
		V_A_CTRL_TT_shadow_intermed_2 <= V_A_CTRL_TT_shadow_intermed_1;
		V_A_CTRL_TT_shadow_intermed_3 <= V_A_CTRL_TT_shadow_intermed_2;
		V_A_CTRL_TT_shadow_intermed_4 <= V_A_CTRL_TT_shadow_intermed_3;
		R_M_CTRL_TT_intermed_1 <= R.M.CTRL.TT;
		RIN_X_CTRL_TT_intermed_1 <= RIN.X.CTRL.TT;
		RIN_X_RESULT6DOWNTO0_intermed_1 <= RIN.X.RESULT ( 6 DOWNTO 0 );
		R_E_CTRL_TT_intermed_1 <= R.E.CTRL.TT;
		R_E_CTRL_TT_intermed_2 <= R_E_CTRL_TT_intermed_1;
		RIN_M_CTRL_TT_intermed_1 <= RIN.M.CTRL.TT;
		RIN_M_CTRL_TT_intermed_2 <= RIN_M_CTRL_TT_intermed_1;
		V_X_RESULT6DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO0_shadow;
		V_M_CTRL_TRAP_shadow_intermed_1 <= V_M_CTRL_TRAP_shadow;
		V_M_CTRL_TRAP_shadow_intermed_2 <= V_M_CTRL_TRAP_shadow_intermed_1;
		RIN_X_CTRL_TRAP_intermed_1 <= RIN.X.CTRL.TRAP;
		V_X_CTRL_TRAP_shadow_intermed_1 <= V_X_CTRL_TRAP_shadow;
		V_A_CTRL_TRAP_shadow_intermed_1 <= V_A_CTRL_TRAP_shadow;
		V_A_CTRL_TRAP_shadow_intermed_2 <= V_A_CTRL_TRAP_shadow_intermed_1;
		V_A_CTRL_TRAP_shadow_intermed_3 <= V_A_CTRL_TRAP_shadow_intermed_2;
		V_A_CTRL_TRAP_shadow_intermed_4 <= V_A_CTRL_TRAP_shadow_intermed_3;
		V_X_MEXC_shadow_intermed_1 <= V_X_MEXC_shadow;
		V_D_MEXC_shadow_intermed_1 <= V_D_MEXC_shadow;
		V_D_MEXC_shadow_intermed_2 <= V_D_MEXC_shadow_intermed_1;
		V_D_MEXC_shadow_intermed_3 <= V_D_MEXC_shadow_intermed_2;
		V_D_MEXC_shadow_intermed_4 <= V_D_MEXC_shadow_intermed_3;
		V_D_MEXC_shadow_intermed_5 <= V_D_MEXC_shadow_intermed_4;
		R_A_CTRL_TRAP_intermed_1 <= R.A.CTRL.TRAP;
		R_A_CTRL_TRAP_intermed_2 <= R_A_CTRL_TRAP_intermed_1;
		R_A_CTRL_TRAP_intermed_3 <= R_A_CTRL_TRAP_intermed_2;
		RIN_X_MEXC_intermed_1 <= RIN.X.MEXC;
		RIN_M_CTRL_TRAP_intermed_1 <= RIN.M.CTRL.TRAP;
		RIN_M_CTRL_TRAP_intermed_2 <= RIN_M_CTRL_TRAP_intermed_1;
		R_M_CTRL_TRAP_intermed_1 <= R.M.CTRL.TRAP;
		ICO_MEXC_intermed_1 <= ICO.MEXC;
		ICO_MEXC_intermed_2 <= ICO_MEXC_intermed_1;
		ICO_MEXC_intermed_3 <= ICO_MEXC_intermed_2;
		ICO_MEXC_intermed_4 <= ICO_MEXC_intermed_3;
		ICO_MEXC_intermed_5 <= ICO_MEXC_intermed_4;
		R_E_CTRL_TRAP_intermed_1 <= R.E.CTRL.TRAP;
		R_E_CTRL_TRAP_intermed_2 <= R_E_CTRL_TRAP_intermed_1;
		RIN_A_CTRL_TRAP_intermed_1 <= RIN.A.CTRL.TRAP;
		RIN_A_CTRL_TRAP_intermed_2 <= RIN_A_CTRL_TRAP_intermed_1;
		RIN_A_CTRL_TRAP_intermed_3 <= RIN_A_CTRL_TRAP_intermed_2;
		RIN_A_CTRL_TRAP_intermed_4 <= RIN_A_CTRL_TRAP_intermed_3;
		V_E_CTRL_TRAP_shadow_intermed_1 <= V_E_CTRL_TRAP_shadow;
		V_E_CTRL_TRAP_shadow_intermed_2 <= V_E_CTRL_TRAP_shadow_intermed_1;
		V_E_CTRL_TRAP_shadow_intermed_3 <= V_E_CTRL_TRAP_shadow_intermed_2;
		RIN_E_CTRL_TRAP_intermed_1 <= RIN.E.CTRL.TRAP;
		RIN_E_CTRL_TRAP_intermed_2 <= RIN_E_CTRL_TRAP_intermed_1;
		RIN_E_CTRL_TRAP_intermed_3 <= RIN_E_CTRL_TRAP_intermed_2;
		RIN_D_MEXC_intermed_1 <= RIN.D.MEXC;
		RIN_D_MEXC_intermed_2 <= RIN_D_MEXC_intermed_1;
		RIN_D_MEXC_intermed_3 <= RIN_D_MEXC_intermed_2;
		RIN_D_MEXC_intermed_4 <= RIN_D_MEXC_intermed_3;
		RIN_D_MEXC_intermed_5 <= RIN_D_MEXC_intermed_4;
		R_D_MEXC_intermed_1 <= R.D.MEXC;
		R_D_MEXC_intermed_2 <= R_D_MEXC_intermed_1;
		R_D_MEXC_intermed_3 <= R_D_MEXC_intermed_2;
		R_D_MEXC_intermed_4 <= R_D_MEXC_intermed_3;
		DCO_MEXC_intermed_1 <= DCO.MEXC;
		DE_INST19_shadow_intermed_1 <= DE_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		V_E_CTRL_INST19_shadow_intermed_1 <= V_E_CTRL_INST19_shadow;
		V_E_CTRL_INST19_shadow_intermed_1 <= V_E_CTRL_INST19_shadow;
		V_E_CTRL_INST19_shadow_intermed_2 <= V_E_CTRL_INST19_shadow_intermed_1;
		R_E_CTRL_INST19_intermed_1 <= R.E.CTRL.INST( 19 );
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST ( 19 );
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST( 19 );
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST ( 19 );
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST( 19 );
		RIN_E_CTRL_INST19_intermed_2 <= RIN_E_CTRL_INST19_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		VP_ERROR_shadow_intermed_1 <= VP_ERROR_shadow;
		RPIN_PWD_intermed_1 <= RPIN.PWD;
		V_X_DEBUG_shadow_intermed_1 <= V_X_DEBUG_shadow;
		VP_PWD_shadow_intermed_1 <= VP_PWD_shadow;
		RPIN_ERROR_intermed_1 <= RPIN.ERROR;
		RIN_X_DEBUG_intermed_1 <= RIN.X.DEBUG;
		VP_ERROR_shadow_intermed_1 <= VP_ERROR_shadow;
		RIN_X_NERROR_intermed_1 <= RIN.X.NERROR;
		RPIN_ERROR_intermed_1 <= RPIN.ERROR;
		V_F_PC31DOWNTO4_shadow_intermed_1 <= V_F_PC31DOWNTO4_shadow;
		V_X_CTRL_TT_shadow_intermed_1 <= V_X_CTRL_TT_shadow;
		V_E_CTRL_TT_shadow_intermed_1 <= V_E_CTRL_TT_shadow;
		V_E_CTRL_TT_shadow_intermed_2 <= V_E_CTRL_TT_shadow_intermed_1;
		V_E_CTRL_TT_shadow_intermed_3 <= V_E_CTRL_TT_shadow_intermed_2;
		RIN_A_CTRL_TT_intermed_1 <= RIN.A.CTRL.TT;
		RIN_A_CTRL_TT_intermed_2 <= RIN_A_CTRL_TT_intermed_1;
		RIN_A_CTRL_TT_intermed_3 <= RIN_A_CTRL_TT_intermed_2;
		RIN_A_CTRL_TT_intermed_4 <= RIN_A_CTRL_TT_intermed_3;
		V_X_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO4_shadow;
		V_X_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO4_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO4_shadow_intermed_3 <= V_X_CTRL_PC31DOWNTO4_shadow_intermed_2;
		IR_ADDR31DOWNTO4_intermed_1 <= IR.ADDR( 31 DOWNTO 4 );
		R_A_CTRL_TT_intermed_1 <= R.A.CTRL.TT;
		R_A_CTRL_TT_intermed_2 <= R_A_CTRL_TT_intermed_1;
		R_A_CTRL_TT_intermed_3 <= R_A_CTRL_TT_intermed_2;
		R_M_CTRL_TT_intermed_1 <= R.M.CTRL.TT;
		RIN_F_PC31DOWNTO4_intermed_1 <= RIN.F.PC( 31 DOWNTO 4 );
		VIR_ADDR31DOWNTO4_shadow_intermed_1 <= VIR_ADDR31DOWNTO4_shadow;
		VIR_ADDR31DOWNTO4_shadow_intermed_2 <= VIR_ADDR31DOWNTO4_shadow_intermed_1;
		RIN_X_RESULT6DOWNTO0_intermed_1 <= RIN.X.RESULT ( 6 DOWNTO 0 );
		R_E_CTRL_TT_intermed_1 <= R.E.CTRL.TT;
		R_E_CTRL_TT_intermed_2 <= R_E_CTRL_TT_intermed_1;
		R_A_CTRL_PC31DOWNTO4_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 4 );
		R_A_CTRL_PC31DOWNTO4_intermed_2 <= R_A_CTRL_PC31DOWNTO4_intermed_1;
		R_A_CTRL_PC31DOWNTO4_intermed_3 <= R_A_CTRL_PC31DOWNTO4_intermed_2;
		R_A_CTRL_PC31DOWNTO4_intermed_4 <= R_A_CTRL_PC31DOWNTO4_intermed_3;
		R_A_CTRL_PC31DOWNTO4_intermed_5 <= R_A_CTRL_PC31DOWNTO4_intermed_4;
		RIN_A_CTRL_PC31DOWNTO4_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 4 );
		RIN_A_CTRL_PC31DOWNTO4_intermed_2 <= RIN_A_CTRL_PC31DOWNTO4_intermed_1;
		RIN_A_CTRL_PC31DOWNTO4_intermed_3 <= RIN_A_CTRL_PC31DOWNTO4_intermed_2;
		RIN_A_CTRL_PC31DOWNTO4_intermed_4 <= RIN_A_CTRL_PC31DOWNTO4_intermed_3;
		RIN_A_CTRL_PC31DOWNTO4_intermed_5 <= RIN_A_CTRL_PC31DOWNTO4_intermed_4;
		RIN_A_CTRL_PC31DOWNTO4_intermed_6 <= RIN_A_CTRL_PC31DOWNTO4_intermed_5;
		R_D_PC31DOWNTO4_intermed_1 <= R.D.PC( 31 DOWNTO 4 );
		R_D_PC31DOWNTO4_intermed_2 <= R_D_PC31DOWNTO4_intermed_1;
		R_D_PC31DOWNTO4_intermed_3 <= R_D_PC31DOWNTO4_intermed_2;
		R_D_PC31DOWNTO4_intermed_4 <= R_D_PC31DOWNTO4_intermed_3;
		R_D_PC31DOWNTO4_intermed_5 <= R_D_PC31DOWNTO4_intermed_4;
		R_D_PC31DOWNTO4_intermed_6 <= R_D_PC31DOWNTO4_intermed_5;
		RIN_X_CTRL_PC31DOWNTO4_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 4 );
		RIN_X_CTRL_PC31DOWNTO4_intermed_2 <= RIN_X_CTRL_PC31DOWNTO4_intermed_1;
		RIN_X_CTRL_PC31DOWNTO4_intermed_3 <= RIN_X_CTRL_PC31DOWNTO4_intermed_2;
		EX_ADD_RES32DOWNTO332DOWNTO5_shadow_intermed_1 <= EX_ADD_RES32DOWNTO332DOWNTO5_shadow;
		V_W_S_TBA_shadow_intermed_1 <= V_W_S_TBA_shadow;
		RIN_M_CTRL_TT_intermed_1 <= RIN.M.CTRL.TT;
		RIN_M_CTRL_TT_intermed_2 <= RIN_M_CTRL_TT_intermed_1;
		RIN_M_CTRL_PC31DOWNTO4_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 4 );
		RIN_M_CTRL_PC31DOWNTO4_intermed_2 <= RIN_M_CTRL_PC31DOWNTO4_intermed_1;
		RIN_M_CTRL_PC31DOWNTO4_intermed_3 <= RIN_M_CTRL_PC31DOWNTO4_intermed_2;
		RIN_M_CTRL_PC31DOWNTO4_intermed_4 <= RIN_M_CTRL_PC31DOWNTO4_intermed_3;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO4_shadow;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO4_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO4_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO4_shadow_intermed_3;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_5 <= V_E_CTRL_PC31DOWNTO4_shadow_intermed_4;
		V_D_PC31DOWNTO4_shadow_intermed_1 <= V_D_PC31DOWNTO4_shadow;
		V_D_PC31DOWNTO4_shadow_intermed_2 <= V_D_PC31DOWNTO4_shadow_intermed_1;
		V_D_PC31DOWNTO4_shadow_intermed_3 <= V_D_PC31DOWNTO4_shadow_intermed_2;
		V_D_PC31DOWNTO4_shadow_intermed_4 <= V_D_PC31DOWNTO4_shadow_intermed_3;
		V_D_PC31DOWNTO4_shadow_intermed_5 <= V_D_PC31DOWNTO4_shadow_intermed_4;
		V_D_PC31DOWNTO4_shadow_intermed_6 <= V_D_PC31DOWNTO4_shadow_intermed_5;
		V_D_PC31DOWNTO4_shadow_intermed_7 <= V_D_PC31DOWNTO4_shadow_intermed_6;
		V_X_RESULT6DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO0_shadow;
		R_X_CTRL_PC31DOWNTO4_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 4 );
		R_X_CTRL_PC31DOWNTO4_intermed_2 <= R_X_CTRL_PC31DOWNTO4_intermed_1;
		V_X_RESULT6DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO0_shadow;
		V_X_RESULT6DOWNTO0_shadow_intermed_2 <= V_X_RESULT6DOWNTO0_shadow_intermed_1;
		RIN_X_RESULT6DOWNTO0_intermed_1 <= RIN.X.RESULT( 6 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO0_intermed_2 <= RIN_X_RESULT6DOWNTO0_intermed_1;
		RIN_E_CTRL_TT_intermed_1 <= RIN.E.CTRL.TT;
		RIN_E_CTRL_TT_intermed_2 <= RIN_E_CTRL_TT_intermed_1;
		RIN_E_CTRL_TT_intermed_3 <= RIN_E_CTRL_TT_intermed_2;
		R_X_RESULT6DOWNTO0_intermed_1 <= R.X.RESULT( 6 DOWNTO 0 );
		V_M_CTRL_TT_shadow_intermed_1 <= V_M_CTRL_TT_shadow;
		V_M_CTRL_TT_shadow_intermed_2 <= V_M_CTRL_TT_shadow_intermed_1;
		IRIN_ADDR31DOWNTO4_intermed_1 <= IRIN.ADDR( 31 DOWNTO 4 );
		IRIN_ADDR31DOWNTO4_intermed_2 <= IRIN_ADDR31DOWNTO4_intermed_1;
		V_M_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO4_shadow;
		V_M_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO4_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO4_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO4_shadow_intermed_2;
		V_M_CTRL_PC31DOWNTO4_shadow_intermed_4 <= V_M_CTRL_PC31DOWNTO4_shadow_intermed_3;
		V_A_CTRL_TT_shadow_intermed_1 <= V_A_CTRL_TT_shadow;
		V_A_CTRL_TT_shadow_intermed_2 <= V_A_CTRL_TT_shadow_intermed_1;
		V_A_CTRL_TT_shadow_intermed_3 <= V_A_CTRL_TT_shadow_intermed_2;
		V_A_CTRL_TT_shadow_intermed_4 <= V_A_CTRL_TT_shadow_intermed_3;
		XC_TRAP_ADDRESS31DOWNTO4_shadow_intermed_1 <= XC_TRAP_ADDRESS31DOWNTO4_shadow;
		R_M_CTRL_PC31DOWNTO4_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 4 );
		R_M_CTRL_PC31DOWNTO4_intermed_2 <= R_M_CTRL_PC31DOWNTO4_intermed_1;
		R_M_CTRL_PC31DOWNTO4_intermed_3 <= R_M_CTRL_PC31DOWNTO4_intermed_2;
		RIN_X_CTRL_TT_intermed_1 <= RIN.X.CTRL.TT;
		RIN_D_PC31DOWNTO4_intermed_1 <= RIN.D.PC( 31 DOWNTO 4 );
		RIN_D_PC31DOWNTO4_intermed_2 <= RIN_D_PC31DOWNTO4_intermed_1;
		RIN_D_PC31DOWNTO4_intermed_3 <= RIN_D_PC31DOWNTO4_intermed_2;
		RIN_D_PC31DOWNTO4_intermed_4 <= RIN_D_PC31DOWNTO4_intermed_3;
		RIN_D_PC31DOWNTO4_intermed_5 <= RIN_D_PC31DOWNTO4_intermed_4;
		RIN_D_PC31DOWNTO4_intermed_6 <= RIN_D_PC31DOWNTO4_intermed_5;
		RIN_D_PC31DOWNTO4_intermed_7 <= RIN_D_PC31DOWNTO4_intermed_6;
		RIN_E_CTRL_PC31DOWNTO4_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 4 );
		RIN_E_CTRL_PC31DOWNTO4_intermed_2 <= RIN_E_CTRL_PC31DOWNTO4_intermed_1;
		RIN_E_CTRL_PC31DOWNTO4_intermed_3 <= RIN_E_CTRL_PC31DOWNTO4_intermed_2;
		RIN_E_CTRL_PC31DOWNTO4_intermed_4 <= RIN_E_CTRL_PC31DOWNTO4_intermed_3;
		RIN_E_CTRL_PC31DOWNTO4_intermed_5 <= RIN_E_CTRL_PC31DOWNTO4_intermed_4;
		EX_JUMP_ADDRESS31DOWNTO4_shadow_intermed_1 <= EX_JUMP_ADDRESS31DOWNTO4_shadow;
		RIN_W_S_TBA_intermed_1 <= RIN.W.S.TBA;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO4_shadow;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_4;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_6 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_5;
		R_E_CTRL_PC31DOWNTO4_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 4 );
		R_E_CTRL_PC31DOWNTO4_intermed_2 <= R_E_CTRL_PC31DOWNTO4_intermed_1;
		R_E_CTRL_PC31DOWNTO4_intermed_3 <= R_E_CTRL_PC31DOWNTO4_intermed_2;
		R_E_CTRL_PC31DOWNTO4_intermed_4 <= R_E_CTRL_PC31DOWNTO4_intermed_3;
		R_D_PC3DOWNTO2_intermed_1 <= R.D.PC( 3 DOWNTO 2 );
		R_D_PC3DOWNTO2_intermed_2 <= R_D_PC3DOWNTO2_intermed_1;
		R_D_PC3DOWNTO2_intermed_3 <= R_D_PC3DOWNTO2_intermed_2;
		R_D_PC3DOWNTO2_intermed_4 <= R_D_PC3DOWNTO2_intermed_3;
		R_D_PC3DOWNTO2_intermed_5 <= R_D_PC3DOWNTO2_intermed_4;
		R_D_PC3DOWNTO2_intermed_6 <= R_D_PC3DOWNTO2_intermed_5;
		V_D_PC3DOWNTO2_shadow_intermed_1 <= V_D_PC3DOWNTO2_shadow;
		V_D_PC3DOWNTO2_shadow_intermed_2 <= V_D_PC3DOWNTO2_shadow_intermed_1;
		V_D_PC3DOWNTO2_shadow_intermed_3 <= V_D_PC3DOWNTO2_shadow_intermed_2;
		V_D_PC3DOWNTO2_shadow_intermed_4 <= V_D_PC3DOWNTO2_shadow_intermed_3;
		V_D_PC3DOWNTO2_shadow_intermed_5 <= V_D_PC3DOWNTO2_shadow_intermed_4;
		V_D_PC3DOWNTO2_shadow_intermed_6 <= V_D_PC3DOWNTO2_shadow_intermed_5;
		V_D_PC3DOWNTO2_shadow_intermed_7 <= V_D_PC3DOWNTO2_shadow_intermed_6;
		VIR_ADDR3DOWNTO2_shadow_intermed_1 <= VIR_ADDR3DOWNTO2_shadow;
		VIR_ADDR3DOWNTO2_shadow_intermed_2 <= VIR_ADDR3DOWNTO2_shadow_intermed_1;
		RIN_D_PC3DOWNTO2_intermed_1 <= RIN.D.PC( 3 DOWNTO 2 );
		RIN_D_PC3DOWNTO2_intermed_2 <= RIN_D_PC3DOWNTO2_intermed_1;
		RIN_D_PC3DOWNTO2_intermed_3 <= RIN_D_PC3DOWNTO2_intermed_2;
		RIN_D_PC3DOWNTO2_intermed_4 <= RIN_D_PC3DOWNTO2_intermed_3;
		RIN_D_PC3DOWNTO2_intermed_5 <= RIN_D_PC3DOWNTO2_intermed_4;
		RIN_D_PC3DOWNTO2_intermed_6 <= RIN_D_PC3DOWNTO2_intermed_5;
		RIN_D_PC3DOWNTO2_intermed_7 <= RIN_D_PC3DOWNTO2_intermed_6;
		R_M_CTRL_PC3DOWNTO2_intermed_1 <= R.M.CTRL.PC( 3 DOWNTO 2 );
		R_M_CTRL_PC3DOWNTO2_intermed_2 <= R_M_CTRL_PC3DOWNTO2_intermed_1;
		R_M_CTRL_PC3DOWNTO2_intermed_3 <= R_M_CTRL_PC3DOWNTO2_intermed_2;
		R_E_CTRL_PC3DOWNTO2_intermed_1 <= R.E.CTRL.PC( 3 DOWNTO 2 );
		R_E_CTRL_PC3DOWNTO2_intermed_2 <= R_E_CTRL_PC3DOWNTO2_intermed_1;
		R_E_CTRL_PC3DOWNTO2_intermed_3 <= R_E_CTRL_PC3DOWNTO2_intermed_2;
		R_E_CTRL_PC3DOWNTO2_intermed_4 <= R_E_CTRL_PC3DOWNTO2_intermed_3;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC3DOWNTO2_shadow;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC3DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC3DOWNTO2_shadow_intermed_2;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_4 <= V_E_CTRL_PC3DOWNTO2_shadow_intermed_3;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_5 <= V_E_CTRL_PC3DOWNTO2_shadow_intermed_4;
		RIN_X_CTRL_PC3DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 3 DOWNTO 2 );
		RIN_X_CTRL_PC3DOWNTO2_intermed_2 <= RIN_X_CTRL_PC3DOWNTO2_intermed_1;
		RIN_X_CTRL_PC3DOWNTO2_intermed_3 <= RIN_X_CTRL_PC3DOWNTO2_intermed_2;
		R_A_CTRL_PC3DOWNTO2_intermed_1 <= R.A.CTRL.PC( 3 DOWNTO 2 );
		R_A_CTRL_PC3DOWNTO2_intermed_2 <= R_A_CTRL_PC3DOWNTO2_intermed_1;
		R_A_CTRL_PC3DOWNTO2_intermed_3 <= R_A_CTRL_PC3DOWNTO2_intermed_2;
		R_A_CTRL_PC3DOWNTO2_intermed_4 <= R_A_CTRL_PC3DOWNTO2_intermed_3;
		R_A_CTRL_PC3DOWNTO2_intermed_5 <= R_A_CTRL_PC3DOWNTO2_intermed_4;
		V_X_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC3DOWNTO2_shadow;
		V_X_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_X_CTRL_PC3DOWNTO2_shadow_intermed_1;
		V_X_CTRL_PC3DOWNTO2_shadow_intermed_3 <= V_X_CTRL_PC3DOWNTO2_shadow_intermed_2;
		RIN_M_CTRL_PC3DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 3 DOWNTO 2 );
		RIN_M_CTRL_PC3DOWNTO2_intermed_2 <= RIN_M_CTRL_PC3DOWNTO2_intermed_1;
		RIN_M_CTRL_PC3DOWNTO2_intermed_3 <= RIN_M_CTRL_PC3DOWNTO2_intermed_2;
		RIN_M_CTRL_PC3DOWNTO2_intermed_4 <= RIN_M_CTRL_PC3DOWNTO2_intermed_3;
		IRIN_ADDR3DOWNTO2_intermed_1 <= IRIN.ADDR( 3 DOWNTO 2 );
		IRIN_ADDR3DOWNTO2_intermed_2 <= IRIN_ADDR3DOWNTO2_intermed_1;
		EX_JUMP_ADDRESS3DOWNTO2_shadow_intermed_1 <= EX_JUMP_ADDRESS3DOWNTO2_shadow;
		EX_ADD_RES32DOWNTO34DOWNTO3_shadow_intermed_1 <= EX_ADD_RES32DOWNTO34DOWNTO3_shadow;
		RIN_A_CTRL_PC3DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 3 DOWNTO 2 );
		RIN_A_CTRL_PC3DOWNTO2_intermed_2 <= RIN_A_CTRL_PC3DOWNTO2_intermed_1;
		RIN_A_CTRL_PC3DOWNTO2_intermed_3 <= RIN_A_CTRL_PC3DOWNTO2_intermed_2;
		RIN_A_CTRL_PC3DOWNTO2_intermed_4 <= RIN_A_CTRL_PC3DOWNTO2_intermed_3;
		RIN_A_CTRL_PC3DOWNTO2_intermed_5 <= RIN_A_CTRL_PC3DOWNTO2_intermed_4;
		RIN_A_CTRL_PC3DOWNTO2_intermed_6 <= RIN_A_CTRL_PC3DOWNTO2_intermed_5;
		XC_TRAP_ADDRESS3DOWNTO2_shadow_intermed_1 <= XC_TRAP_ADDRESS3DOWNTO2_shadow;
		V_F_PC3DOWNTO2_shadow_intermed_1 <= V_F_PC3DOWNTO2_shadow;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC3DOWNTO2_shadow;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_3;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_5 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_4;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_6 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_5;
		IR_ADDR3DOWNTO2_intermed_1 <= IR.ADDR( 3 DOWNTO 2 );
		V_M_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC3DOWNTO2_shadow;
		V_M_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC3DOWNTO2_shadow_intermed_1;
		V_M_CTRL_PC3DOWNTO2_shadow_intermed_3 <= V_M_CTRL_PC3DOWNTO2_shadow_intermed_2;
		V_M_CTRL_PC3DOWNTO2_shadow_intermed_4 <= V_M_CTRL_PC3DOWNTO2_shadow_intermed_3;
		R_X_CTRL_PC3DOWNTO2_intermed_1 <= R.X.CTRL.PC( 3 DOWNTO 2 );
		R_X_CTRL_PC3DOWNTO2_intermed_2 <= R_X_CTRL_PC3DOWNTO2_intermed_1;
		RIN_E_CTRL_PC3DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 3 DOWNTO 2 );
		RIN_E_CTRL_PC3DOWNTO2_intermed_2 <= RIN_E_CTRL_PC3DOWNTO2_intermed_1;
		RIN_E_CTRL_PC3DOWNTO2_intermed_3 <= RIN_E_CTRL_PC3DOWNTO2_intermed_2;
		RIN_E_CTRL_PC3DOWNTO2_intermed_4 <= RIN_E_CTRL_PC3DOWNTO2_intermed_3;
		RIN_E_CTRL_PC3DOWNTO2_intermed_5 <= RIN_E_CTRL_PC3DOWNTO2_intermed_4;
		RIN_F_PC3DOWNTO2_intermed_1 <= RIN.F.PC( 3 DOWNTO 2 );
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_X_DEBUG_intermed_1 <= RIN.X.DEBUG;
		RIN_D_PC_intermed_1 <= RIN.D.PC;
		RIN_D_PC_intermed_2 <= RIN_D_PC_intermed_1;
		RIN_D_PC_intermed_3 <= RIN_D_PC_intermed_2;
		RIN_D_PC_intermed_4 <= RIN_D_PC_intermed_3;
		RIN_D_PC_intermed_5 <= RIN_D_PC_intermed_4;
		RIN_A_CTRL_PC_intermed_1 <= RIN.A.CTRL.PC;
		RIN_A_CTRL_PC_intermed_2 <= RIN_A_CTRL_PC_intermed_1;
		RIN_A_CTRL_PC_intermed_3 <= RIN_A_CTRL_PC_intermed_2;
		RIN_A_CTRL_PC_intermed_4 <= RIN_A_CTRL_PC_intermed_3;
		R_A_CTRL_PC_intermed_1 <= R.A.CTRL.PC;
		R_A_CTRL_PC_intermed_2 <= R_A_CTRL_PC_intermed_1;
		R_A_CTRL_PC_intermed_3 <= R_A_CTRL_PC_intermed_2;
		V_E_CTRL_PC_shadow_intermed_1 <= V_E_CTRL_PC_shadow;
		V_E_CTRL_PC_shadow_intermed_2 <= V_E_CTRL_PC_shadow_intermed_1;
		V_E_CTRL_PC_shadow_intermed_3 <= V_E_CTRL_PC_shadow_intermed_2;
		R_M_CTRL_PC_intermed_1 <= R.M.CTRL.PC;
		R_E_CTRL_PC_intermed_1 <= R.E.CTRL.PC;
		R_E_CTRL_PC_intermed_2 <= R_E_CTRL_PC_intermed_1;
		RIN_M_CTRL_PC_intermed_1 <= RIN.M.CTRL.PC;
		RIN_M_CTRL_PC_intermed_2 <= RIN_M_CTRL_PC_intermed_1;
		V_X_CTRL_PC_shadow_intermed_1 <= V_X_CTRL_PC_shadow;
		V_M_CTRL_PC_shadow_intermed_1 <= V_M_CTRL_PC_shadow;
		V_M_CTRL_PC_shadow_intermed_2 <= V_M_CTRL_PC_shadow_intermed_1;
		V_A_CTRL_PC_shadow_intermed_1 <= V_A_CTRL_PC_shadow;
		V_A_CTRL_PC_shadow_intermed_2 <= V_A_CTRL_PC_shadow_intermed_1;
		V_A_CTRL_PC_shadow_intermed_3 <= V_A_CTRL_PC_shadow_intermed_2;
		V_A_CTRL_PC_shadow_intermed_4 <= V_A_CTRL_PC_shadow_intermed_3;
		R_D_PC_intermed_1 <= R.D.PC;
		R_D_PC_intermed_2 <= R_D_PC_intermed_1;
		R_D_PC_intermed_3 <= R_D_PC_intermed_2;
		R_D_PC_intermed_4 <= R_D_PC_intermed_3;
		RIN_E_CTRL_PC_intermed_1 <= RIN.E.CTRL.PC;
		RIN_E_CTRL_PC_intermed_2 <= RIN_E_CTRL_PC_intermed_1;
		RIN_E_CTRL_PC_intermed_3 <= RIN_E_CTRL_PC_intermed_2;
		RIN_X_CTRL_PC_intermed_1 <= RIN.X.CTRL.PC;
		V_D_PC_shadow_intermed_1 <= V_D_PC_shadow;
		V_D_PC_shadow_intermed_2 <= V_D_PC_shadow_intermed_1;
		V_D_PC_shadow_intermed_3 <= V_D_PC_shadow_intermed_2;
		V_D_PC_shadow_intermed_4 <= V_D_PC_shadow_intermed_3;
		V_D_PC_shadow_intermed_5 <= V_D_PC_shadow_intermed_4;
		IRIN_ADDR_intermed_1 <= IRIN.ADDR;
		V_E_CTRL_TT_shadow_intermed_1 <= V_E_CTRL_TT_shadow;
		V_E_CTRL_TT_shadow_intermed_2 <= V_E_CTRL_TT_shadow_intermed_1;
		V_E_CTRL_TT_shadow_intermed_3 <= V_E_CTRL_TT_shadow_intermed_2;
		V_X_CTRL_TT_shadow_intermed_1 <= V_X_CTRL_TT_shadow;
		RIN_A_CTRL_TT_intermed_1 <= RIN.A.CTRL.TT;
		RIN_A_CTRL_TT_intermed_2 <= RIN_A_CTRL_TT_intermed_1;
		RIN_A_CTRL_TT_intermed_3 <= RIN_A_CTRL_TT_intermed_2;
		RIN_A_CTRL_TT_intermed_4 <= RIN_A_CTRL_TT_intermed_3;
		R_A_CTRL_TT_intermed_1 <= R.A.CTRL.TT;
		R_A_CTRL_TT_intermed_2 <= R_A_CTRL_TT_intermed_1;
		R_A_CTRL_TT_intermed_3 <= R_A_CTRL_TT_intermed_2;
		R_M_CTRL_TT_intermed_1 <= R.M.CTRL.TT;
		RIN_X_RESULT6DOWNTO0_intermed_1 <= RIN.X.RESULT ( 6 DOWNTO 0 );
		DSUIN_TT_intermed_1 <= DSUIN.TT;
		R_E_CTRL_TT_intermed_1 <= R.E.CTRL.TT;
		R_E_CTRL_TT_intermed_2 <= R_E_CTRL_TT_intermed_1;
		RIN_M_CTRL_TT_intermed_1 <= RIN.M.CTRL.TT;
		RIN_M_CTRL_TT_intermed_2 <= RIN_M_CTRL_TT_intermed_1;
		V_X_RESULT6DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO0_shadow;
		V_X_RESULT6DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO0_shadow;
		V_X_RESULT6DOWNTO0_shadow_intermed_2 <= V_X_RESULT6DOWNTO0_shadow_intermed_1;
		RIN_X_RESULT6DOWNTO0_intermed_1 <= RIN.X.RESULT( 6 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO0_intermed_2 <= RIN_X_RESULT6DOWNTO0_intermed_1;
		RIN_E_CTRL_TT_intermed_1 <= RIN.E.CTRL.TT;
		RIN_E_CTRL_TT_intermed_2 <= RIN_E_CTRL_TT_intermed_1;
		RIN_E_CTRL_TT_intermed_3 <= RIN_E_CTRL_TT_intermed_2;
		V_M_CTRL_TT_shadow_intermed_1 <= V_M_CTRL_TT_shadow;
		V_M_CTRL_TT_shadow_intermed_2 <= V_M_CTRL_TT_shadow_intermed_1;
		R_X_RESULT6DOWNTO0_intermed_1 <= R.X.RESULT( 6 DOWNTO 0 );
		V_A_CTRL_TT_shadow_intermed_1 <= V_A_CTRL_TT_shadow;
		V_A_CTRL_TT_shadow_intermed_2 <= V_A_CTRL_TT_shadow_intermed_1;
		V_A_CTRL_TT_shadow_intermed_3 <= V_A_CTRL_TT_shadow_intermed_2;
		V_A_CTRL_TT_shadow_intermed_4 <= V_A_CTRL_TT_shadow_intermed_3;
		RIN_X_CTRL_TT_intermed_1 <= RIN.X.CTRL.TT;
		RPIN_PWD_intermed_1 <= RPIN.PWD;
		IRIN_PWD_intermed_1 <= IRIN.PWD;
		V_E_CTRL_TT_shadow_intermed_1 <= V_E_CTRL_TT_shadow;
		V_E_CTRL_TT_shadow_intermed_2 <= V_E_CTRL_TT_shadow_intermed_1;
		V_E_CTRL_TT_shadow_intermed_3 <= V_E_CTRL_TT_shadow_intermed_2;
		V_X_CTRL_TT_shadow_intermed_1 <= V_X_CTRL_TT_shadow;
		RIN_A_CTRL_TT_intermed_1 <= RIN.A.CTRL.TT;
		RIN_A_CTRL_TT_intermed_2 <= RIN_A_CTRL_TT_intermed_1;
		RIN_A_CTRL_TT_intermed_3 <= RIN_A_CTRL_TT_intermed_2;
		RIN_A_CTRL_TT_intermed_4 <= RIN_A_CTRL_TT_intermed_3;
		R_A_CTRL_TT_intermed_1 <= R.A.CTRL.TT;
		R_A_CTRL_TT_intermed_2 <= R_A_CTRL_TT_intermed_1;
		R_A_CTRL_TT_intermed_3 <= R_A_CTRL_TT_intermed_2;
		R_M_CTRL_TT_intermed_1 <= R.M.CTRL.TT;
		RIN_X_RESULT6DOWNTO0_intermed_1 <= RIN.X.RESULT ( 6 DOWNTO 0 );
		R_E_CTRL_TT_intermed_1 <= R.E.CTRL.TT;
		R_E_CTRL_TT_intermed_2 <= R_E_CTRL_TT_intermed_1;
		RIN_M_CTRL_TT_intermed_1 <= RIN.M.CTRL.TT;
		RIN_M_CTRL_TT_intermed_2 <= RIN_M_CTRL_TT_intermed_1;
		V_X_RESULT6DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO0_shadow;
		V_X_RESULT6DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO0_shadow;
		V_X_RESULT6DOWNTO0_shadow_intermed_2 <= V_X_RESULT6DOWNTO0_shadow_intermed_1;
		RIN_X_RESULT6DOWNTO0_intermed_1 <= RIN.X.RESULT( 6 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO0_intermed_2 <= RIN_X_RESULT6DOWNTO0_intermed_1;
		RIN_E_CTRL_TT_intermed_1 <= RIN.E.CTRL.TT;
		RIN_E_CTRL_TT_intermed_2 <= RIN_E_CTRL_TT_intermed_1;
		RIN_E_CTRL_TT_intermed_3 <= RIN_E_CTRL_TT_intermed_2;
		V_M_CTRL_TT_shadow_intermed_1 <= V_M_CTRL_TT_shadow;
		V_M_CTRL_TT_shadow_intermed_2 <= V_M_CTRL_TT_shadow_intermed_1;
		R_X_RESULT6DOWNTO0_intermed_1 <= R.X.RESULT( 6 DOWNTO 0 );
		RIN_W_S_TT_intermed_1 <= RIN.W.S.TT;
		V_A_CTRL_TT_shadow_intermed_1 <= V_A_CTRL_TT_shadow;
		V_A_CTRL_TT_shadow_intermed_2 <= V_A_CTRL_TT_shadow_intermed_1;
		V_A_CTRL_TT_shadow_intermed_3 <= V_A_CTRL_TT_shadow_intermed_2;
		V_A_CTRL_TT_shadow_intermed_4 <= V_A_CTRL_TT_shadow_intermed_3;
		RIN_X_CTRL_TT_intermed_1 <= RIN.X.CTRL.TT;
		RIN_W_S_S_intermed_1 <= RIN.W.S.S;
		RIN_W_S_PS_intermed_1 <= RIN.W.S.PS;
		V_W_S_S_shadow_intermed_1 <= V_W_S_S_shadow;
		RIN_W_S_S_intermed_1 <= RIN.W.S.S;
		RIN_E_CTRL_RD6DOWNTO0_intermed_1 <= RIN.E.CTRL.RD( 6 DOWNTO 0 );
		RIN_E_CTRL_RD6DOWNTO0_intermed_2 <= RIN_E_CTRL_RD6DOWNTO0_intermed_1;
		RIN_E_CTRL_RD6DOWNTO0_intermed_3 <= RIN_E_CTRL_RD6DOWNTO0_intermed_2;
		RIN_M_CTRL_RD6DOWNTO0_intermed_1 <= RIN.M.CTRL.RD( 6 DOWNTO 0 );
		RIN_M_CTRL_RD6DOWNTO0_intermed_2 <= RIN_M_CTRL_RD6DOWNTO0_intermed_1;
		RIN_X_CTRL_RD6DOWNTO0_intermed_1 <= RIN.X.CTRL.RD( 6 DOWNTO 0 );
		V_X_CTRL_RD6DOWNTO0_shadow_intermed_1 <= V_X_CTRL_RD6DOWNTO0_shadow;
		RIN_W_S_CWP_intermed_1 <= RIN.W.S.CWP;
		V_M_CTRL_RD6DOWNTO0_shadow_intermed_1 <= V_M_CTRL_RD6DOWNTO0_shadow;
		V_M_CTRL_RD6DOWNTO0_shadow_intermed_2 <= V_M_CTRL_RD6DOWNTO0_shadow_intermed_1;
		R_E_CTRL_RD6DOWNTO0_intermed_1 <= R.E.CTRL.RD( 6 DOWNTO 0 );
		R_E_CTRL_RD6DOWNTO0_intermed_2 <= R_E_CTRL_RD6DOWNTO0_intermed_1;
		V_E_CTRL_RD6DOWNTO0_shadow_intermed_1 <= V_E_CTRL_RD6DOWNTO0_shadow;
		V_E_CTRL_RD6DOWNTO0_shadow_intermed_2 <= V_E_CTRL_RD6DOWNTO0_shadow_intermed_1;
		V_E_CTRL_RD6DOWNTO0_shadow_intermed_3 <= V_E_CTRL_RD6DOWNTO0_shadow_intermed_2;
		V_A_CTRL_RD6DOWNTO0_shadow_intermed_1 <= V_A_CTRL_RD6DOWNTO0_shadow;
		V_A_CTRL_RD6DOWNTO0_shadow_intermed_2 <= V_A_CTRL_RD6DOWNTO0_shadow_intermed_1;
		V_A_CTRL_RD6DOWNTO0_shadow_intermed_3 <= V_A_CTRL_RD6DOWNTO0_shadow_intermed_2;
		V_A_CTRL_RD6DOWNTO0_shadow_intermed_4 <= V_A_CTRL_RD6DOWNTO0_shadow_intermed_3;
		R_A_CTRL_RD6DOWNTO0_intermed_1 <= R.A.CTRL.RD( 6 DOWNTO 0 );
		R_A_CTRL_RD6DOWNTO0_intermed_2 <= R_A_CTRL_RD6DOWNTO0_intermed_1;
		R_A_CTRL_RD6DOWNTO0_intermed_3 <= R_A_CTRL_RD6DOWNTO0_intermed_2;
		RIN_A_CTRL_RD6DOWNTO0_intermed_1 <= RIN.A.CTRL.RD( 6 DOWNTO 0 );
		RIN_A_CTRL_RD6DOWNTO0_intermed_2 <= RIN_A_CTRL_RD6DOWNTO0_intermed_1;
		RIN_A_CTRL_RD6DOWNTO0_intermed_3 <= RIN_A_CTRL_RD6DOWNTO0_intermed_2;
		RIN_A_CTRL_RD6DOWNTO0_intermed_4 <= RIN_A_CTRL_RD6DOWNTO0_intermed_3;
		R_M_CTRL_RD6DOWNTO0_intermed_1 <= R.M.CTRL.RD( 6 DOWNTO 0 );
		V_W_S_CWP_shadow_intermed_1 <= V_W_S_CWP_shadow;
		RIN_W_S_ET_intermed_1 <= RIN.W.S.ET;
		RIN_W_S_CWP_intermed_1 <= RIN.W.S.CWP;
		RPIN_ERROR_intermed_1 <= RPIN.ERROR;
		RIN_D_PC_intermed_1 <= RIN.D.PC;
		RIN_D_PC_intermed_2 <= RIN_D_PC_intermed_1;
		RIN_D_PC_intermed_3 <= RIN_D_PC_intermed_2;
		RIN_D_PC_intermed_4 <= RIN_D_PC_intermed_3;
		RIN_D_PC_intermed_5 <= RIN_D_PC_intermed_4;
		RIN_D_PC_intermed_6 <= RIN_D_PC_intermed_5;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_3 <= RIN_M_CTRL_PC31DOWNTO2_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_4 <= RIN_M_CTRL_PC31DOWNTO2_intermed_3;
		VIR_ADDR_shadow_intermed_1 <= VIR_ADDR_shadow;
		RIN_A_CTRL_PC_intermed_1 <= RIN.A.CTRL.PC;
		RIN_A_CTRL_PC_intermed_2 <= RIN_A_CTRL_PC_intermed_1;
		RIN_A_CTRL_PC_intermed_3 <= RIN_A_CTRL_PC_intermed_2;
		RIN_A_CTRL_PC_intermed_4 <= RIN_A_CTRL_PC_intermed_3;
		RIN_A_CTRL_PC_intermed_5 <= RIN_A_CTRL_PC_intermed_4;
		R_A_CTRL_PC_intermed_1 <= R.A.CTRL.PC;
		R_A_CTRL_PC_intermed_2 <= R_A_CTRL_PC_intermed_1;
		R_A_CTRL_PC_intermed_3 <= R_A_CTRL_PC_intermed_2;
		R_A_CTRL_PC_intermed_4 <= R_A_CTRL_PC_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_5 <= V_D_PC31DOWNTO2_shadow_intermed_4;
		V_D_PC31DOWNTO2_shadow_intermed_6 <= V_D_PC31DOWNTO2_shadow_intermed_5;
		V_D_PC31DOWNTO2_shadow_intermed_7 <= V_D_PC31DOWNTO2_shadow_intermed_6;
		V_E_CTRL_PC_shadow_intermed_1 <= V_E_CTRL_PC_shadow;
		V_E_CTRL_PC_shadow_intermed_2 <= V_E_CTRL_PC_shadow_intermed_1;
		V_E_CTRL_PC_shadow_intermed_3 <= V_E_CTRL_PC_shadow_intermed_2;
		V_E_CTRL_PC_shadow_intermed_4 <= V_E_CTRL_PC_shadow_intermed_3;
		EX_ADD_RES32DOWNTO3_shadow_intermed_1 <= EX_ADD_RES32DOWNTO3_shadow;
		XC_TRAP_ADDRESS_shadow_intermed_1 <= XC_TRAP_ADDRESS_shadow;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_5 <= RIN_D_PC31DOWNTO2_intermed_4;
		RIN_D_PC31DOWNTO2_intermed_6 <= RIN_D_PC31DOWNTO2_intermed_5;
		RIN_D_PC31DOWNTO2_intermed_7 <= RIN_D_PC31DOWNTO2_intermed_6;
		EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_1 <= EX_ADD_RES32DOWNTO332DOWNTO3_shadow;
		V_F_PC31DOWNTO2_shadow_intermed_1 <= V_F_PC31DOWNTO2_shadow;
		RIN_F_PC31DOWNTO2_intermed_1 <= RIN.F.PC( 31 DOWNTO 2 );
		R_M_CTRL_PC_intermed_1 <= R.M.CTRL.PC;
		R_M_CTRL_PC_intermed_2 <= R_M_CTRL_PC_intermed_1;
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_2 <= RIN_X_CTRL_PC31DOWNTO2_intermed_1;
		RIN_X_CTRL_PC31DOWNTO2_intermed_3 <= RIN_X_CTRL_PC31DOWNTO2_intermed_2;
		R_X_CTRL_PC_intermed_1 <= R.X.CTRL.PC;
		R_E_CTRL_PC_intermed_1 <= R.E.CTRL.PC;
		R_E_CTRL_PC_intermed_2 <= R_E_CTRL_PC_intermed_1;
		R_E_CTRL_PC_intermed_3 <= R_E_CTRL_PC_intermed_2;
		IRIN_ADDR31DOWNTO2_intermed_1 <= IRIN.ADDR( 31 DOWNTO 2 );
		IRIN_ADDR31DOWNTO2_intermed_2 <= IRIN_ADDR31DOWNTO2_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_6 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_5;
		RIN_M_CTRL_PC_intermed_1 <= RIN.M.CTRL.PC;
		RIN_M_CTRL_PC_intermed_2 <= RIN_M_CTRL_PC_intermed_1;
		RIN_M_CTRL_PC_intermed_3 <= RIN_M_CTRL_PC_intermed_2;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		R_D_PC31DOWNTO2_intermed_4 <= R_D_PC31DOWNTO2_intermed_3;
		R_D_PC31DOWNTO2_intermed_5 <= R_D_PC31DOWNTO2_intermed_4;
		R_D_PC31DOWNTO2_intermed_6 <= R_D_PC31DOWNTO2_intermed_5;
		VIR_ADDR31DOWNTO2_shadow_intermed_1 <= VIR_ADDR31DOWNTO2_shadow;
		VIR_ADDR31DOWNTO2_shadow_intermed_2 <= VIR_ADDR31DOWNTO2_shadow_intermed_1;
		V_X_CTRL_PC_shadow_intermed_1 <= V_X_CTRL_PC_shadow;
		V_X_CTRL_PC_shadow_intermed_2 <= V_X_CTRL_PC_shadow_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 2 );
		R_M_CTRL_PC31DOWNTO2_intermed_2 <= R_M_CTRL_PC31DOWNTO2_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_3 <= R_M_CTRL_PC31DOWNTO2_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_4;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		RIN_A_CTRL_PC31DOWNTO2_intermed_5 <= RIN_A_CTRL_PC31DOWNTO2_intermed_4;
		RIN_A_CTRL_PC31DOWNTO2_intermed_6 <= RIN_A_CTRL_PC31DOWNTO2_intermed_5;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_4 <= R_A_CTRL_PC31DOWNTO2_intermed_3;
		R_A_CTRL_PC31DOWNTO2_intermed_5 <= R_A_CTRL_PC31DOWNTO2_intermed_4;
		V_M_CTRL_PC_shadow_intermed_1 <= V_M_CTRL_PC_shadow;
		V_M_CTRL_PC_shadow_intermed_2 <= V_M_CTRL_PC_shadow_intermed_1;
		V_M_CTRL_PC_shadow_intermed_3 <= V_M_CTRL_PC_shadow_intermed_2;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_A_CTRL_PC_shadow_intermed_1 <= V_A_CTRL_PC_shadow;
		V_A_CTRL_PC_shadow_intermed_2 <= V_A_CTRL_PC_shadow_intermed_1;
		V_A_CTRL_PC_shadow_intermed_3 <= V_A_CTRL_PC_shadow_intermed_2;
		V_A_CTRL_PC_shadow_intermed_4 <= V_A_CTRL_PC_shadow_intermed_3;
		V_A_CTRL_PC_shadow_intermed_5 <= V_A_CTRL_PC_shadow_intermed_4;
		R_X_CTRL_PC31DOWNTO2_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 2 );
		R_X_CTRL_PC31DOWNTO2_intermed_2 <= R_X_CTRL_PC31DOWNTO2_intermed_1;
		R_D_PC_intermed_1 <= R.D.PC;
		R_D_PC_intermed_2 <= R_D_PC_intermed_1;
		R_D_PC_intermed_3 <= R_D_PC_intermed_2;
		R_D_PC_intermed_4 <= R_D_PC_intermed_3;
		R_D_PC_intermed_5 <= R_D_PC_intermed_4;
		RIN_F_PC_intermed_1 <= RIN.F.PC;
		XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_1 <= XC_TRAP_ADDRESS31DOWNTO2_shadow;
		RIN_E_CTRL_PC_intermed_1 <= RIN.E.CTRL.PC;
		RIN_E_CTRL_PC_intermed_2 <= RIN_E_CTRL_PC_intermed_1;
		RIN_E_CTRL_PC_intermed_3 <= RIN_E_CTRL_PC_intermed_2;
		RIN_E_CTRL_PC_intermed_4 <= RIN_E_CTRL_PC_intermed_3;
		RIN_X_CTRL_PC_intermed_1 <= RIN.X.CTRL.PC;
		RIN_X_CTRL_PC_intermed_2 <= RIN_X_CTRL_PC_intermed_1;
		V_D_PC_shadow_intermed_1 <= V_D_PC_shadow;
		V_D_PC_shadow_intermed_2 <= V_D_PC_shadow_intermed_1;
		V_D_PC_shadow_intermed_3 <= V_D_PC_shadow_intermed_2;
		V_D_PC_shadow_intermed_4 <= V_D_PC_shadow_intermed_3;
		V_D_PC_shadow_intermed_5 <= V_D_PC_shadow_intermed_4;
		V_D_PC_shadow_intermed_6 <= V_D_PC_shadow_intermed_5;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_3 <= R_E_CTRL_PC31DOWNTO2_intermed_2;
		R_E_CTRL_PC31DOWNTO2_intermed_4 <= R_E_CTRL_PC31DOWNTO2_intermed_3;
		IRIN_ADDR_intermed_1 <= IRIN.ADDR;
		EX_JUMP_ADDRESS_shadow_intermed_1 <= EX_JUMP_ADDRESS_shadow;
		EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_1 <= EX_JUMP_ADDRESS31DOWNTO2_shadow;
		IR_ADDR31DOWNTO2_intermed_1 <= IR.ADDR( 31 DOWNTO 2 );
		V_F_PC_shadow_intermed_1 <= V_F_PC_shadow;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_4 <= RIN_E_CTRL_PC31DOWNTO2_intermed_3;
		RIN_E_CTRL_PC31DOWNTO2_intermed_5 <= RIN_E_CTRL_PC31DOWNTO2_intermed_4;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO2_shadow;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_2;
		DSUIN_TBUFCNT_intermed_1 <= DSUIN.TBUFCNT;
		RIN_W_EXCEPT_intermed_1 <= RIN.W.EXCEPT;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_3 <= RIN_M_CTRL_PC31DOWNTO2_intermed_2;
		RIN_X_RESULT_intermed_1 <= RIN.X.RESULT;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO2_shadow;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC ( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_5 <= V_D_PC31DOWNTO2_shadow_intermed_4;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_5 <= RIN_D_PC31DOWNTO2_intermed_4;
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC ( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC ( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC ( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_2 <= RIN_X_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC ( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		R_D_PC31DOWNTO2_intermed_4 <= R_D_PC31DOWNTO2_intermed_3;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC ( 31 DOWNTO 2 );
		DCO_DATA0_intermed_1 <= DCO.DATA ( 0 );
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		V_X_DATA0_shadow_intermed_2 <= V_X_DATA0_shadow_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 2 );
		R_M_CTRL_PC31DOWNTO2_intermed_2 <= R_M_CTRL_PC31DOWNTO2_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		RIN_A_CTRL_PC31DOWNTO2_intermed_5 <= RIN_A_CTRL_PC31DOWNTO2_intermed_4;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_4 <= R_A_CTRL_PC31DOWNTO2_intermed_3;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2;
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA ( 0 );
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC ( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		V_X_RESULT_shadow_intermed_1 <= V_X_RESULT_shadow;
		R_X_CTRL_PC31DOWNTO2_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 2 );
		RIN_W_RESULT_intermed_1 <= RIN.W.RESULT;
		R_X_DATA0_intermed_1 <= R.X.DATA( 0 );
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_3 <= R_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_4 <= RIN_E_CTRL_PC31DOWNTO2_intermed_3;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO2_shadow;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA( 0 );
		RIN_X_DATA0_intermed_2 <= RIN_X_DATA0_intermed_1;
		V_M_CTRL_RD7DOWNTO0_shadow_intermed_1 <= V_M_CTRL_RD7DOWNTO0_shadow;
		V_M_CTRL_RD7DOWNTO0_shadow_intermed_2 <= V_M_CTRL_RD7DOWNTO0_shadow_intermed_1;
		V_E_CTRL_RD7DOWNTO0_shadow_intermed_1 <= V_E_CTRL_RD7DOWNTO0_shadow;
		V_E_CTRL_RD7DOWNTO0_shadow_intermed_2 <= V_E_CTRL_RD7DOWNTO0_shadow_intermed_1;
		V_E_CTRL_RD7DOWNTO0_shadow_intermed_3 <= V_E_CTRL_RD7DOWNTO0_shadow_intermed_2;
		R_E_CTRL_RD7DOWNTO0_intermed_1 <= R.E.CTRL.RD ( 7 DOWNTO 0 );
		R_E_CTRL_RD7DOWNTO0_intermed_2 <= R_E_CTRL_RD7DOWNTO0_intermed_1;
		V_X_CTRL_RD7DOWNTO0_shadow_intermed_1 <= V_X_CTRL_RD7DOWNTO0_shadow;
		V_A_CTRL_RD7DOWNTO0_shadow_intermed_1 <= V_A_CTRL_RD7DOWNTO0_shadow;
		V_A_CTRL_RD7DOWNTO0_shadow_intermed_2 <= V_A_CTRL_RD7DOWNTO0_shadow_intermed_1;
		V_A_CTRL_RD7DOWNTO0_shadow_intermed_3 <= V_A_CTRL_RD7DOWNTO0_shadow_intermed_2;
		V_A_CTRL_RD7DOWNTO0_shadow_intermed_4 <= V_A_CTRL_RD7DOWNTO0_shadow_intermed_3;
		RIN_W_WA_intermed_1 <= RIN.W.WA;
		RIN_A_CTRL_RD7DOWNTO0_intermed_1 <= RIN.A.CTRL.RD ( 7 DOWNTO 0 );
		RIN_A_CTRL_RD7DOWNTO0_intermed_2 <= RIN_A_CTRL_RD7DOWNTO0_intermed_1;
		RIN_A_CTRL_RD7DOWNTO0_intermed_3 <= RIN_A_CTRL_RD7DOWNTO0_intermed_2;
		RIN_A_CTRL_RD7DOWNTO0_intermed_4 <= RIN_A_CTRL_RD7DOWNTO0_intermed_3;
		R_M_CTRL_RD7DOWNTO0_intermed_1 <= R.M.CTRL.RD ( 7 DOWNTO 0 );
		R_A_CTRL_RD7DOWNTO0_intermed_1 <= R.A.CTRL.RD ( 7 DOWNTO 0 );
		R_A_CTRL_RD7DOWNTO0_intermed_2 <= R_A_CTRL_RD7DOWNTO0_intermed_1;
		R_A_CTRL_RD7DOWNTO0_intermed_3 <= R_A_CTRL_RD7DOWNTO0_intermed_2;
		RIN_E_CTRL_RD7DOWNTO0_intermed_1 <= RIN.E.CTRL.RD ( 7 DOWNTO 0 );
		RIN_E_CTRL_RD7DOWNTO0_intermed_2 <= RIN_E_CTRL_RD7DOWNTO0_intermed_1;
		RIN_E_CTRL_RD7DOWNTO0_intermed_3 <= RIN_E_CTRL_RD7DOWNTO0_intermed_2;
		RIN_X_CTRL_RD7DOWNTO0_intermed_1 <= RIN.X.CTRL.RD ( 7 DOWNTO 0 );
		RIN_M_CTRL_RD7DOWNTO0_intermed_1 <= RIN.M.CTRL.RD ( 7 DOWNTO 0 );
		RIN_M_CTRL_RD7DOWNTO0_intermed_2 <= RIN_M_CTRL_RD7DOWNTO0_intermed_1;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_A_CTRL_ANNUL_intermed_2 <= RIN_A_CTRL_ANNUL_intermed_1;
		RIN_A_CTRL_ANNUL_intermed_3 <= RIN_A_CTRL_ANNUL_intermed_2;
		RIN_A_CTRL_ANNUL_intermed_4 <= RIN_A_CTRL_ANNUL_intermed_3;
		RIN_A_CTRL_ANNUL_intermed_5 <= RIN_A_CTRL_ANNUL_intermed_4;
		R_A_CTRL_ANNUL_intermed_1 <= R.A.CTRL.ANNUL;
		R_A_CTRL_ANNUL_intermed_2 <= R_A_CTRL_ANNUL_intermed_1;
		R_A_CTRL_ANNUL_intermed_3 <= R_A_CTRL_ANNUL_intermed_2;
		R_A_CTRL_ANNUL_intermed_4 <= R_A_CTRL_ANNUL_intermed_3;
		R_X_ANNUL_ALL_intermed_1 <= R.X.ANNUL_ALL;
		R_X_ANNUL_ALL_intermed_2 <= R_X_ANNUL_ALL_intermed_1;
		R_X_ANNUL_ALL_intermed_3 <= R_X_ANNUL_ALL_intermed_2;
		R_X_ANNUL_ALL_intermed_4 <= R_X_ANNUL_ALL_intermed_3;
		V_X_CTRL_WREG_shadow_intermed_1 <= V_X_CTRL_WREG_shadow;
		RIN_X_CTRL_WREG_intermed_1 <= RIN.X.CTRL.WREG;
		RIN_M_CTRL_WREG_intermed_1 <= RIN.M.CTRL.WREG;
		RIN_M_CTRL_WREG_intermed_2 <= RIN_M_CTRL_WREG_intermed_1;
		RIN_A_CTRL_WREG_intermed_1 <= RIN.A.CTRL.WREG;
		RIN_A_CTRL_WREG_intermed_2 <= RIN_A_CTRL_WREG_intermed_1;
		RIN_A_CTRL_WREG_intermed_3 <= RIN_A_CTRL_WREG_intermed_2;
		RIN_A_CTRL_WREG_intermed_4 <= RIN_A_CTRL_WREG_intermed_3;
		V_A_CTRL_WREG_shadow_intermed_1 <= V_A_CTRL_WREG_shadow;
		V_A_CTRL_WREG_shadow_intermed_2 <= V_A_CTRL_WREG_shadow_intermed_1;
		V_A_CTRL_WREG_shadow_intermed_3 <= V_A_CTRL_WREG_shadow_intermed_2;
		V_A_CTRL_WREG_shadow_intermed_4 <= V_A_CTRL_WREG_shadow_intermed_3;
		R_A_CTRL_WREG_intermed_1 <= R.A.CTRL.WREG;
		R_A_CTRL_WREG_intermed_2 <= R_A_CTRL_WREG_intermed_1;
		R_A_CTRL_WREG_intermed_3 <= R_A_CTRL_WREG_intermed_2;
		RIN_W_WREG_intermed_1 <= RIN.W.WREG;
		V_X_ANNUL_ALL_shadow_intermed_1 <= V_X_ANNUL_ALL_shadow;
		V_X_ANNUL_ALL_shadow_intermed_2 <= V_X_ANNUL_ALL_shadow_intermed_1;
		V_X_ANNUL_ALL_shadow_intermed_3 <= V_X_ANNUL_ALL_shadow_intermed_2;
		V_X_ANNUL_ALL_shadow_intermed_4 <= V_X_ANNUL_ALL_shadow_intermed_3;
		R_M_CTRL_WREG_intermed_1 <= R.M.CTRL.WREG;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_X_ANNUL_ALL_intermed_2 <= RIN_X_ANNUL_ALL_intermed_1;
		RIN_X_ANNUL_ALL_intermed_3 <= RIN_X_ANNUL_ALL_intermed_2;
		RIN_X_ANNUL_ALL_intermed_4 <= RIN_X_ANNUL_ALL_intermed_3;
		RIN_X_ANNUL_ALL_intermed_5 <= RIN_X_ANNUL_ALL_intermed_4;
		V_M_CTRL_WREG_shadow_intermed_1 <= V_M_CTRL_WREG_shadow;
		V_M_CTRL_WREG_shadow_intermed_2 <= V_M_CTRL_WREG_shadow_intermed_1;
		R_E_CTRL_WREG_intermed_1 <= R.E.CTRL.WREG;
		R_E_CTRL_WREG_intermed_2 <= R_E_CTRL_WREG_intermed_1;
		V_A_CTRL_ANNUL_shadow_intermed_1 <= V_A_CTRL_ANNUL_shadow;
		V_A_CTRL_ANNUL_shadow_intermed_2 <= V_A_CTRL_ANNUL_shadow_intermed_1;
		V_A_CTRL_ANNUL_shadow_intermed_3 <= V_A_CTRL_ANNUL_shadow_intermed_2;
		V_A_CTRL_ANNUL_shadow_intermed_4 <= V_A_CTRL_ANNUL_shadow_intermed_3;
		RIN_E_CTRL_WREG_intermed_1 <= RIN.E.CTRL.WREG;
		RIN_E_CTRL_WREG_intermed_2 <= RIN_E_CTRL_WREG_intermed_1;
		RIN_E_CTRL_WREG_intermed_3 <= RIN_E_CTRL_WREG_intermed_2;
		V_E_CTRL_WREG_shadow_intermed_1 <= V_E_CTRL_WREG_shadow;
		V_E_CTRL_WREG_shadow_intermed_2 <= V_E_CTRL_WREG_shadow_intermed_1;
		V_E_CTRL_WREG_shadow_intermed_3 <= V_E_CTRL_WREG_shadow_intermed_2;
		RIN_W_S_SVT_intermed_1 <= RIN.W.S.SVT;
		RIN_W_S_DWT_intermed_1 <= RIN.W.S.DWT;
		RIN_W_S_EF_intermed_1 <= RIN.W.S.EF;
		RIN_E_CTRL_intermed_1 <= RIN.E.CTRL;
		RIN_E_CTRL_intermed_2 <= RIN_E_CTRL_intermed_1;
		R_E_CTRL_intermed_1 <= R.E.CTRL;
		RIN_X_CTRL_intermed_1 <= RIN.X.CTRL;
		RIN_M_CTRL_intermed_1 <= RIN.M.CTRL;
		V_E_CTRL_shadow_intermed_1 <= V_E_CTRL_shadow;
		V_E_CTRL_shadow_intermed_2 <= V_E_CTRL_shadow_intermed_1;
		RIN_A_CTRL_intermed_1 <= RIN.A.CTRL;
		RIN_A_CTRL_intermed_2 <= RIN_A_CTRL_intermed_1;
		RIN_A_CTRL_intermed_3 <= RIN_A_CTRL_intermed_2;
		V_M_CTRL_shadow_intermed_1 <= V_M_CTRL_shadow;
		V_A_CTRL_shadow_intermed_1 <= V_A_CTRL_shadow;
		V_A_CTRL_shadow_intermed_2 <= V_A_CTRL_shadow_intermed_1;
		V_A_CTRL_shadow_intermed_3 <= V_A_CTRL_shadow_intermed_2;
		R_A_CTRL_intermed_1 <= R.A.CTRL;
		R_A_CTRL_intermed_2 <= R_A_CTRL_intermed_1;
		V_M_DCI_shadow_intermed_1 <= V_M_DCI_shadow;
		RIN_M_DCI_intermed_1 <= RIN.M.DCI;
		RIN_X_DCI_intermed_1 <= RIN.X.DCI;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_A_CTRL_ANNUL_intermed_2 <= RIN_A_CTRL_ANNUL_intermed_1;
		RIN_A_CTRL_ANNUL_intermed_3 <= RIN_A_CTRL_ANNUL_intermed_2;
		RIN_A_CTRL_ANNUL_intermed_4 <= RIN_A_CTRL_ANNUL_intermed_3;
		R_A_CTRL_ANNUL_intermed_1 <= R.A.CTRL.ANNUL;
		R_A_CTRL_ANNUL_intermed_2 <= R_A_CTRL_ANNUL_intermed_1;
		R_A_CTRL_ANNUL_intermed_3 <= R_A_CTRL_ANNUL_intermed_2;
		RIN_M_CTRL_RETT_intermed_1 <= RIN.M.CTRL.RETT;
		V_M_CTRL_ANNUL_shadow_intermed_1 <= V_M_CTRL_ANNUL_shadow;
		R_X_ANNUL_ALL_intermed_1 <= R.X.ANNUL_ALL;
		R_X_ANNUL_ALL_intermed_2 <= R_X_ANNUL_ALL_intermed_1;
		R_X_ANNUL_ALL_intermed_3 <= R_X_ANNUL_ALL_intermed_2;
		RIN_M_CTRL_ANNUL_intermed_1 <= RIN.M.CTRL.ANNUL;
		V_E_CTRL_RETT_shadow_intermed_1 <= V_E_CTRL_RETT_shadow;
		V_E_CTRL_RETT_shadow_intermed_2 <= V_E_CTRL_RETT_shadow_intermed_1;
		V_A_CTRL_RETT_shadow_intermed_1 <= V_A_CTRL_RETT_shadow;
		V_A_CTRL_RETT_shadow_intermed_2 <= V_A_CTRL_RETT_shadow_intermed_1;
		V_A_CTRL_RETT_shadow_intermed_3 <= V_A_CTRL_RETT_shadow_intermed_2;
		RIN_A_CTRL_RETT_intermed_1 <= RIN.A.CTRL.RETT;
		RIN_A_CTRL_RETT_intermed_2 <= RIN_A_CTRL_RETT_intermed_1;
		RIN_A_CTRL_RETT_intermed_3 <= RIN_A_CTRL_RETT_intermed_2;
		V_X_ANNUL_ALL_shadow_intermed_1 <= V_X_ANNUL_ALL_shadow;
		V_X_ANNUL_ALL_shadow_intermed_2 <= V_X_ANNUL_ALL_shadow_intermed_1;
		V_X_ANNUL_ALL_shadow_intermed_3 <= V_X_ANNUL_ALL_shadow_intermed_2;
		RIN_E_CTRL_ANNUL_intermed_1 <= RIN.E.CTRL.ANNUL;
		RIN_E_CTRL_ANNUL_intermed_2 <= RIN_E_CTRL_ANNUL_intermed_1;
		R_E_CTRL_RETT_intermed_1 <= R.E.CTRL.RETT;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_X_ANNUL_ALL_intermed_2 <= RIN_X_ANNUL_ALL_intermed_1;
		RIN_X_ANNUL_ALL_intermed_3 <= RIN_X_ANNUL_ALL_intermed_2;
		RIN_X_ANNUL_ALL_intermed_4 <= RIN_X_ANNUL_ALL_intermed_3;
		RIN_E_CTRL_RETT_intermed_1 <= RIN.E.CTRL.RETT;
		RIN_E_CTRL_RETT_intermed_2 <= RIN_E_CTRL_RETT_intermed_1;
		V_E_CTRL_ANNUL_shadow_intermed_1 <= V_E_CTRL_ANNUL_shadow;
		V_E_CTRL_ANNUL_shadow_intermed_2 <= V_E_CTRL_ANNUL_shadow_intermed_1;
		V_A_CTRL_ANNUL_shadow_intermed_1 <= V_A_CTRL_ANNUL_shadow;
		V_A_CTRL_ANNUL_shadow_intermed_2 <= V_A_CTRL_ANNUL_shadow_intermed_1;
		V_A_CTRL_ANNUL_shadow_intermed_3 <= V_A_CTRL_ANNUL_shadow_intermed_2;
		RIN_X_CTRL_RETT_intermed_1 <= RIN.X.CTRL.RETT;
		V_M_CTRL_RETT_shadow_intermed_1 <= V_M_CTRL_RETT_shadow;
		R_A_CTRL_RETT_intermed_1 <= R.A.CTRL.RETT;
		R_A_CTRL_RETT_intermed_2 <= R_A_CTRL_RETT_intermed_1;
		R_E_CTRL_ANNUL_intermed_1 <= R.E.CTRL.ANNUL;
		V_E_MAC_shadow_intermed_1 <= V_E_MAC_shadow;
		V_E_MAC_shadow_intermed_2 <= V_E_MAC_shadow_intermed_1;
		RIN_M_MAC_intermed_1 <= RIN.M.MAC;
		RIN_E_MAC_intermed_1 <= RIN.E.MAC;
		RIN_E_MAC_intermed_2 <= RIN_E_MAC_intermed_1;
		R_E_MAC_intermed_1 <= R.E.MAC;
		V_M_MAC_shadow_intermed_1 <= V_M_MAC_shadow;
		RIN_X_MAC_intermed_1 <= RIN.X.MAC;
		V_M_RESULT1DOWNTO0_shadow_intermed_1 <= V_M_RESULT1DOWNTO0_shadow;
		V_M_RESULT1DOWNTO0_shadow_intermed_2 <= V_M_RESULT1DOWNTO0_shadow_intermed_1;
		RIN_X_LADDR_intermed_1 <= RIN.X.LADDR;
		RIN_M_RESULT1DOWNTO0_intermed_1 <= RIN.M.RESULT( 1 DOWNTO 0 );
		RIN_M_RESULT1DOWNTO0_intermed_2 <= RIN_M_RESULT1DOWNTO0_intermed_1;
		V_M_RESULT1DOWNTO0_shadow_intermed_1 <= V_M_RESULT1DOWNTO0_shadow;
		R_M_RESULT1DOWNTO0_intermed_1 <= R.M.RESULT( 1 DOWNTO 0 );
		RIN_M_RESULT1DOWNTO0_intermed_1 <= RIN.M.RESULT ( 1 DOWNTO 0 );
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_A_CTRL_ANNUL_intermed_2 <= RIN_A_CTRL_ANNUL_intermed_1;
		RIN_A_CTRL_ANNUL_intermed_3 <= RIN_A_CTRL_ANNUL_intermed_2;
		R_A_CTRL_ANNUL_intermed_1 <= R.A.CTRL.ANNUL;
		R_A_CTRL_ANNUL_intermed_2 <= R_A_CTRL_ANNUL_intermed_1;
		V_M_CTRL_ANNUL_shadow_intermed_1 <= V_M_CTRL_ANNUL_shadow;
		R_X_ANNUL_ALL_intermed_1 <= R.X.ANNUL_ALL;
		RIN_X_CTRL_ANNUL_intermed_1 <= RIN.X.CTRL.ANNUL;
		RIN_M_CTRL_ANNUL_intermed_1 <= RIN.M.CTRL.ANNUL;
		V_X_ANNUL_ALL_shadow_intermed_1 <= V_X_ANNUL_ALL_shadow;
		RIN_E_CTRL_ANNUL_intermed_1 <= RIN.E.CTRL.ANNUL;
		RIN_E_CTRL_ANNUL_intermed_2 <= RIN_E_CTRL_ANNUL_intermed_1;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_X_ANNUL_ALL_intermed_2 <= RIN_X_ANNUL_ALL_intermed_1;
		V_E_CTRL_ANNUL_shadow_intermed_1 <= V_E_CTRL_ANNUL_shadow;
		V_E_CTRL_ANNUL_shadow_intermed_2 <= V_E_CTRL_ANNUL_shadow_intermed_1;
		V_A_CTRL_ANNUL_shadow_intermed_1 <= V_A_CTRL_ANNUL_shadow;
		V_A_CTRL_ANNUL_shadow_intermed_2 <= V_A_CTRL_ANNUL_shadow_intermed_1;
		V_A_CTRL_ANNUL_shadow_intermed_3 <= V_A_CTRL_ANNUL_shadow_intermed_2;
		R_E_CTRL_ANNUL_intermed_1 <= R.E.CTRL.ANNUL;
		V_E_CTRL_TT_shadow_intermed_1 <= V_E_CTRL_TT_shadow;
		V_E_CTRL_TT_shadow_intermed_2 <= V_E_CTRL_TT_shadow_intermed_1;
		V_E_CTRL_TT_shadow_intermed_3 <= V_E_CTRL_TT_shadow_intermed_2;
		RIN_A_CTRL_TT_intermed_1 <= RIN.A.CTRL.TT;
		RIN_A_CTRL_TT_intermed_2 <= RIN_A_CTRL_TT_intermed_1;
		RIN_A_CTRL_TT_intermed_3 <= RIN_A_CTRL_TT_intermed_2;
		RIN_A_CTRL_TT_intermed_4 <= RIN_A_CTRL_TT_intermed_3;
		R_A_CTRL_TT_intermed_1 <= R.A.CTRL.TT;
		R_A_CTRL_TT_intermed_2 <= R_A_CTRL_TT_intermed_1;
		R_A_CTRL_TT_intermed_3 <= R_A_CTRL_TT_intermed_2;
		R_M_CTRL_TT_intermed_1 <= R.M.CTRL.TT;
		R_E_CTRL_TT_intermed_1 <= R.E.CTRL.TT;
		R_E_CTRL_TT_intermed_2 <= R_E_CTRL_TT_intermed_1;
		RIN_M_CTRL_TT_intermed_1 <= RIN.M.CTRL.TT;
		RIN_M_CTRL_TT_intermed_2 <= RIN_M_CTRL_TT_intermed_1;
		RIN_E_CTRL_TT_intermed_1 <= RIN.E.CTRL.TT;
		RIN_E_CTRL_TT_intermed_2 <= RIN_E_CTRL_TT_intermed_1;
		RIN_E_CTRL_TT_intermed_3 <= RIN_E_CTRL_TT_intermed_2;
		V_M_CTRL_TT_shadow_intermed_1 <= V_M_CTRL_TT_shadow;
		V_M_CTRL_TT_shadow_intermed_2 <= V_M_CTRL_TT_shadow_intermed_1;
		V_A_CTRL_TT_shadow_intermed_1 <= V_A_CTRL_TT_shadow;
		V_A_CTRL_TT_shadow_intermed_2 <= V_A_CTRL_TT_shadow_intermed_1;
		V_A_CTRL_TT_shadow_intermed_3 <= V_A_CTRL_TT_shadow_intermed_2;
		V_A_CTRL_TT_shadow_intermed_4 <= V_A_CTRL_TT_shadow_intermed_3;
		RIN_X_CTRL_TT_intermed_1 <= RIN.X.CTRL.TT;
		V_X_DATA0_shadow_intermed_1 <= V_X_DATA0_shadow;
		V_X_DATA0_shadow_intermed_2 <= V_X_DATA0_shadow_intermed_1;
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA ( 0 );
		R_X_DATA0_intermed_1 <= R.X.DATA( 0 );
		RIN_X_DATA0_intermed_1 <= RIN.X.DATA( 0 );
		RIN_X_DATA0_intermed_2 <= RIN_X_DATA0_intermed_1;
		V_X_DATA1_shadow_intermed_1 <= V_X_DATA1_shadow;
		V_X_DATA1_shadow_intermed_2 <= V_X_DATA1_shadow_intermed_1;
		RIN_X_DATA1_intermed_1 <= RIN.X.DATA ( 1 );
		R_X_DATA1_intermed_1 <= R.X.DATA( 1 );
		RIN_X_DATA1_intermed_1 <= RIN.X.DATA( 1 );
		RIN_X_DATA1_intermed_2 <= RIN_X_DATA1_intermed_1;
		RIN_X_SET_intermed_1 <= RIN.X.SET;
		V_M_DCI_SIZE_shadow_intermed_1 <= V_M_DCI_SIZE_shadow;
		V_M_DCI_SIZE_shadow_intermed_2 <= V_M_DCI_SIZE_shadow_intermed_1;
		R_M_DCI_SIZE_intermed_1 <= R.M.DCI.SIZE;
		RIN_X_DCI_SIZE_intermed_1 <= RIN.X.DCI.SIZE;
		RIN_M_DCI_SIZE_intermed_1 <= RIN.M.DCI.SIZE;
		RIN_M_DCI_SIZE_intermed_2 <= RIN_M_DCI_SIZE_intermed_1;
		RIN_M_DCI_SIGNED_intermed_1 <= RIN.M.DCI.SIGNED;
		RIN_M_DCI_SIGNED_intermed_2 <= RIN_M_DCI_SIGNED_intermed_1;
		R_M_DCI_SIGNED_intermed_1 <= R.M.DCI.SIGNED;
		RIN_X_DCI_SIGNED_intermed_1 <= RIN.X.DCI.SIGNED;
		V_M_DCI_SIGNED_shadow_intermed_1 <= V_M_DCI_SIGNED_shadow;
		V_M_DCI_SIGNED_shadow_intermed_2 <= V_M_DCI_SIGNED_shadow_intermed_1;
		RIN_X_MEXC_intermed_1 <= RIN.X.MEXC;
		RIN_X_ICC_intermed_1 <= RIN.X.ICC;
		R_A_CTRL_WICC_intermed_1 <= R.A.CTRL.WICC;
		R_A_CTRL_WICC_intermed_2 <= R_A_CTRL_WICC_intermed_1;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_A_CTRL_ANNUL_intermed_2 <= RIN_A_CTRL_ANNUL_intermed_1;
		RIN_A_CTRL_ANNUL_intermed_3 <= RIN_A_CTRL_ANNUL_intermed_2;
		RIN_A_CTRL_ANNUL_intermed_4 <= RIN_A_CTRL_ANNUL_intermed_3;
		V_E_CTRL_WICC_shadow_intermed_1 <= V_E_CTRL_WICC_shadow;
		V_E_CTRL_WICC_shadow_intermed_2 <= V_E_CTRL_WICC_shadow_intermed_1;
		V_A_CTRL_WICC_shadow_intermed_1 <= V_A_CTRL_WICC_shadow;
		V_A_CTRL_WICC_shadow_intermed_2 <= V_A_CTRL_WICC_shadow_intermed_1;
		V_A_CTRL_WICC_shadow_intermed_3 <= V_A_CTRL_WICC_shadow_intermed_2;
		R_A_CTRL_ANNUL_intermed_1 <= R.A.CTRL.ANNUL;
		R_A_CTRL_ANNUL_intermed_2 <= R_A_CTRL_ANNUL_intermed_1;
		R_A_CTRL_ANNUL_intermed_3 <= R_A_CTRL_ANNUL_intermed_2;
		RIN_X_CTRL_WICC_intermed_1 <= RIN.X.CTRL.WICC;
		R_X_ANNUL_ALL_intermed_1 <= R.X.ANNUL_ALL;
		R_X_ANNUL_ALL_intermed_2 <= R_X_ANNUL_ALL_intermed_1;
		R_X_ANNUL_ALL_intermed_3 <= R_X_ANNUL_ALL_intermed_2;
		RIN_E_CTRL_WICC_intermed_1 <= RIN.E.CTRL.WICC;
		RIN_E_CTRL_WICC_intermed_2 <= RIN_E_CTRL_WICC_intermed_1;
		RIN_M_CTRL_WICC_intermed_1 <= RIN.M.CTRL.WICC;
		R_E_CTRL_WICC_intermed_1 <= R.E.CTRL.WICC;
		V_X_ANNUL_ALL_shadow_intermed_1 <= V_X_ANNUL_ALL_shadow;
		V_X_ANNUL_ALL_shadow_intermed_2 <= V_X_ANNUL_ALL_shadow_intermed_1;
		V_X_ANNUL_ALL_shadow_intermed_3 <= V_X_ANNUL_ALL_shadow_intermed_2;
		V_M_CTRL_WICC_shadow_intermed_1 <= V_M_CTRL_WICC_shadow;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_X_ANNUL_ALL_intermed_2 <= RIN_X_ANNUL_ALL_intermed_1;
		RIN_X_ANNUL_ALL_intermed_3 <= RIN_X_ANNUL_ALL_intermed_2;
		RIN_X_ANNUL_ALL_intermed_4 <= RIN_X_ANNUL_ALL_intermed_3;
		RIN_A_CTRL_WICC_intermed_1 <= RIN.A.CTRL.WICC;
		RIN_A_CTRL_WICC_intermed_2 <= RIN_A_CTRL_WICC_intermed_1;
		RIN_A_CTRL_WICC_intermed_3 <= RIN_A_CTRL_WICC_intermed_2;
		V_A_CTRL_ANNUL_shadow_intermed_1 <= V_A_CTRL_ANNUL_shadow;
		V_A_CTRL_ANNUL_shadow_intermed_2 <= V_A_CTRL_ANNUL_shadow_intermed_1;
		V_A_CTRL_ANNUL_shadow_intermed_3 <= V_A_CTRL_ANNUL_shadow_intermed_2;
		RIN_E_CTRL_intermed_1 <= RIN.E.CTRL;
		RIN_M_CTRL_intermed_1 <= RIN.M.CTRL;
		V_E_CTRL_shadow_intermed_1 <= V_E_CTRL_shadow;
		RIN_A_CTRL_intermed_1 <= RIN.A.CTRL;
		RIN_A_CTRL_intermed_2 <= RIN_A_CTRL_intermed_1;
		V_A_CTRL_shadow_intermed_1 <= V_A_CTRL_shadow;
		V_A_CTRL_shadow_intermed_2 <= V_A_CTRL_shadow_intermed_1;
		R_A_CTRL_intermed_1 <= R.A.CTRL;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_A_CTRL_ANNUL_intermed_2 <= RIN_A_CTRL_ANNUL_intermed_1;
		RIN_A_CTRL_ANNUL_intermed_3 <= RIN_A_CTRL_ANNUL_intermed_2;
		R_A_CTRL_ANNUL_intermed_1 <= R.A.CTRL.ANNUL;
		R_A_CTRL_ANNUL_intermed_2 <= R_A_CTRL_ANNUL_intermed_1;
		RIN_M_CTRL_RETT_intermed_1 <= RIN.M.CTRL.RETT;
		R_X_ANNUL_ALL_intermed_1 <= R.X.ANNUL_ALL;
		R_X_ANNUL_ALL_intermed_2 <= R_X_ANNUL_ALL_intermed_1;
		V_E_CTRL_RETT_shadow_intermed_1 <= V_E_CTRL_RETT_shadow;
		V_A_CTRL_RETT_shadow_intermed_1 <= V_A_CTRL_RETT_shadow;
		V_A_CTRL_RETT_shadow_intermed_2 <= V_A_CTRL_RETT_shadow_intermed_1;
		RIN_A_CTRL_RETT_intermed_1 <= RIN.A.CTRL.RETT;
		RIN_A_CTRL_RETT_intermed_2 <= RIN_A_CTRL_RETT_intermed_1;
		V_X_ANNUL_ALL_shadow_intermed_1 <= V_X_ANNUL_ALL_shadow;
		V_X_ANNUL_ALL_shadow_intermed_2 <= V_X_ANNUL_ALL_shadow_intermed_1;
		RIN_E_CTRL_ANNUL_intermed_1 <= RIN.E.CTRL.ANNUL;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_X_ANNUL_ALL_intermed_2 <= RIN_X_ANNUL_ALL_intermed_1;
		RIN_X_ANNUL_ALL_intermed_3 <= RIN_X_ANNUL_ALL_intermed_2;
		RIN_E_CTRL_RETT_intermed_1 <= RIN.E.CTRL.RETT;
		V_E_CTRL_ANNUL_shadow_intermed_1 <= V_E_CTRL_ANNUL_shadow;
		V_A_CTRL_ANNUL_shadow_intermed_1 <= V_A_CTRL_ANNUL_shadow;
		V_A_CTRL_ANNUL_shadow_intermed_2 <= V_A_CTRL_ANNUL_shadow_intermed_1;
		R_A_CTRL_RETT_intermed_1 <= R.A.CTRL.RETT;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_A_CTRL_ANNUL_intermed_2 <= RIN_A_CTRL_ANNUL_intermed_1;
		RIN_A_CTRL_ANNUL_intermed_3 <= RIN_A_CTRL_ANNUL_intermed_2;
		R_A_CTRL_ANNUL_intermed_1 <= R.A.CTRL.ANNUL;
		R_A_CTRL_ANNUL_intermed_2 <= R_A_CTRL_ANNUL_intermed_1;
		R_X_ANNUL_ALL_intermed_1 <= R.X.ANNUL_ALL;
		R_X_ANNUL_ALL_intermed_2 <= R_X_ANNUL_ALL_intermed_1;
		RIN_M_CTRL_WREG_intermed_1 <= RIN.M.CTRL.WREG;
		RIN_A_CTRL_WREG_intermed_1 <= RIN.A.CTRL.WREG;
		RIN_A_CTRL_WREG_intermed_2 <= RIN_A_CTRL_WREG_intermed_1;
		V_A_CTRL_WREG_shadow_intermed_1 <= V_A_CTRL_WREG_shadow;
		V_A_CTRL_WREG_shadow_intermed_2 <= V_A_CTRL_WREG_shadow_intermed_1;
		R_A_CTRL_WREG_intermed_1 <= R.A.CTRL.WREG;
		V_X_ANNUL_ALL_shadow_intermed_1 <= V_X_ANNUL_ALL_shadow;
		V_X_ANNUL_ALL_shadow_intermed_2 <= V_X_ANNUL_ALL_shadow_intermed_1;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_X_ANNUL_ALL_intermed_2 <= RIN_X_ANNUL_ALL_intermed_1;
		RIN_X_ANNUL_ALL_intermed_3 <= RIN_X_ANNUL_ALL_intermed_2;
		V_A_CTRL_ANNUL_shadow_intermed_1 <= V_A_CTRL_ANNUL_shadow;
		V_A_CTRL_ANNUL_shadow_intermed_2 <= V_A_CTRL_ANNUL_shadow_intermed_1;
		RIN_E_CTRL_WREG_intermed_1 <= RIN.E.CTRL.WREG;
		V_E_CTRL_WREG_shadow_intermed_1 <= V_E_CTRL_WREG_shadow;
		RIN_E_CWP_intermed_1 <= RIN.E.CWP;
		V_A_CWP_shadow_intermed_1 <= V_A_CWP_shadow;
		RIN_D_CWP_intermed_1 <= RIN.D.CWP;
		RIN_D_CWP_intermed_2 <= RIN_D_CWP_intermed_1;
		RIN_A_CWP_intermed_1 <= RIN.A.CWP;
		V_D_CWP_shadow_intermed_1 <= V_D_CWP_shadow;
		V_D_CWP_shadow_intermed_2 <= V_D_CWP_shadow_intermed_1;
		R_D_CWP_intermed_1 <= R.D.CWP;
		R_A_SU_intermed_1 <= R.A.SU;
		RIN_A_SU_intermed_1 <= RIN.A.SU;
		RIN_A_SU_intermed_2 <= RIN_A_SU_intermed_1;
		V_E_SU_shadow_intermed_1 <= V_E_SU_shadow;
		V_A_SU_shadow_intermed_1 <= V_A_SU_shadow;
		V_A_SU_shadow_intermed_2 <= V_A_SU_shadow_intermed_1;
		RIN_M_SU_intermed_1 <= RIN.M.SU;
		RIN_E_SU_intermed_1 <= RIN.E.SU;
		RIN_M_MUL_intermed_1 <= RIN.M.MUL;
		RIN_M_NALIGN_intermed_1 <= RIN.M.NALIGN;
		V_X_DATA03_shadow_intermed_1 <= V_X_DATA03_shadow;
		V_X_DATA03_shadow_intermed_2 <= V_X_DATA03_shadow_intermed_1;
		V_X_DATA03_shadow_intermed_1 <= V_X_DATA03_shadow;
		DCO_DATA03_intermed_1 <= DCO.DATA ( 0 )( 3 );
		RIN_X_DATA03_intermed_1 <= RIN.X.DATA ( 0 )( 3 );
		R_X_DATA03_intermed_1 <= R.X.DATA( 0 )( 3 );
		RIN_X_DATA03_intermed_1 <= RIN.X.DATA( 0 )( 3 );
		RIN_X_DATA03_intermed_2 <= RIN_X_DATA03_intermed_1;
		RIN_E_OP23_intermed_1 <= RIN.E.OP2( 3 );
		RIN_E_OP13_intermed_1 <= RIN.E.OP1( 3 );
		V_E_OP23_shadow_intermed_1 <= V_E_OP23_shadow;
		V_E_OP13_shadow_intermed_1 <= V_E_OP13_shadow;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_A_CTRL_ANNUL_intermed_2 <= RIN_A_CTRL_ANNUL_intermed_1;
		RIN_A_CTRL_ANNUL_intermed_3 <= RIN_A_CTRL_ANNUL_intermed_2;
		R_A_CTRL_ANNUL_intermed_1 <= R.A.CTRL.ANNUL;
		R_A_CTRL_ANNUL_intermed_2 <= R_A_CTRL_ANNUL_intermed_1;
		RIN_M_CTRL_ANNUL_intermed_1 <= RIN.M.CTRL.ANNUL;
		RIN_E_CTRL_ANNUL_intermed_1 <= RIN.E.CTRL.ANNUL;
		RIN_E_CTRL_ANNUL_intermed_2 <= RIN_E_CTRL_ANNUL_intermed_1;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		V_E_CTRL_ANNUL_shadow_intermed_1 <= V_E_CTRL_ANNUL_shadow;
		V_E_CTRL_ANNUL_shadow_intermed_2 <= V_E_CTRL_ANNUL_shadow_intermed_1;
		V_A_CTRL_ANNUL_shadow_intermed_1 <= V_A_CTRL_ANNUL_shadow;
		V_A_CTRL_ANNUL_shadow_intermed_2 <= V_A_CTRL_ANNUL_shadow_intermed_1;
		V_A_CTRL_ANNUL_shadow_intermed_3 <= V_A_CTRL_ANNUL_shadow_intermed_2;
		R_E_CTRL_ANNUL_intermed_1 <= R.E.CTRL.ANNUL;
		R_A_CTRL_WICC_intermed_1 <= R.A.CTRL.WICC;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_A_CTRL_ANNUL_intermed_2 <= RIN_A_CTRL_ANNUL_intermed_1;
		RIN_A_CTRL_ANNUL_intermed_3 <= RIN_A_CTRL_ANNUL_intermed_2;
		V_E_CTRL_WICC_shadow_intermed_1 <= V_E_CTRL_WICC_shadow;
		V_A_CTRL_WICC_shadow_intermed_1 <= V_A_CTRL_WICC_shadow;
		V_A_CTRL_WICC_shadow_intermed_2 <= V_A_CTRL_WICC_shadow_intermed_1;
		R_A_CTRL_ANNUL_intermed_1 <= R.A.CTRL.ANNUL;
		R_A_CTRL_ANNUL_intermed_2 <= R_A_CTRL_ANNUL_intermed_1;
		R_X_ANNUL_ALL_intermed_1 <= R.X.ANNUL_ALL;
		R_X_ANNUL_ALL_intermed_2 <= R_X_ANNUL_ALL_intermed_1;
		RIN_E_CTRL_WICC_intermed_1 <= RIN.E.CTRL.WICC;
		RIN_M_CTRL_WICC_intermed_1 <= RIN.M.CTRL.WICC;
		V_X_ANNUL_ALL_shadow_intermed_1 <= V_X_ANNUL_ALL_shadow;
		V_X_ANNUL_ALL_shadow_intermed_2 <= V_X_ANNUL_ALL_shadow_intermed_1;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_X_ANNUL_ALL_intermed_2 <= RIN_X_ANNUL_ALL_intermed_1;
		RIN_X_ANNUL_ALL_intermed_3 <= RIN_X_ANNUL_ALL_intermed_2;
		RIN_A_CTRL_WICC_intermed_1 <= RIN.A.CTRL.WICC;
		RIN_A_CTRL_WICC_intermed_2 <= RIN_A_CTRL_WICC_intermed_1;
		V_A_CTRL_ANNUL_shadow_intermed_1 <= V_A_CTRL_ANNUL_shadow;
		V_A_CTRL_ANNUL_shadow_intermed_2 <= V_A_CTRL_ANNUL_shadow_intermed_1;
		V_E_MAC_shadow_intermed_1 <= V_E_MAC_shadow;
		RIN_M_MAC_intermed_1 <= RIN.M.MAC;
		RIN_E_MAC_intermed_1 <= RIN.E.MAC;
		R_A_CTRL_LD_intermed_1 <= R.A.CTRL.LD;
		R_A_CTRL_LD_intermed_2 <= R_A_CTRL_LD_intermed_1;
		RIN_A_CTRL_LD_intermed_1 <= RIN.A.CTRL.LD;
		RIN_A_CTRL_LD_intermed_2 <= RIN_A_CTRL_LD_intermed_1;
		RIN_A_CTRL_LD_intermed_3 <= RIN_A_CTRL_LD_intermed_2;
		V_E_CTRL_LD_shadow_intermed_1 <= V_E_CTRL_LD_shadow;
		V_E_CTRL_LD_shadow_intermed_2 <= V_E_CTRL_LD_shadow_intermed_1;
		R_E_CTRL_LD_intermed_1 <= R.E.CTRL.LD;
		RIN_E_CTRL_LD_intermed_1 <= RIN.E.CTRL.LD;
		RIN_E_CTRL_LD_intermed_2 <= RIN_E_CTRL_LD_intermed_1;
		RIN_M_CTRL_LD_intermed_1 <= RIN.M.CTRL.LD;
		V_A_CTRL_LD_shadow_intermed_1 <= V_A_CTRL_LD_shadow;
		V_A_CTRL_LD_shadow_intermed_2 <= V_A_CTRL_LD_shadow_intermed_1;
		V_A_CTRL_LD_shadow_intermed_3 <= V_A_CTRL_LD_shadow_intermed_2;
		RIN_E_CTRL_intermed_1 <= RIN.E.CTRL;
		RIN_A_CTRL_intermed_1 <= RIN.A.CTRL;
		V_A_CTRL_shadow_intermed_1 <= V_A_CTRL_shadow;
		RIN_E_JMPL_intermed_1 <= RIN.E.JMPL;
		RIN_A_JMPL_intermed_1 <= RIN.A.JMPL;
		V_A_JMPL_shadow_intermed_1 <= V_A_JMPL_shadow;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		R_X_ANNUL_ALL_intermed_1 <= R.X.ANNUL_ALL;
		V_X_ANNUL_ALL_shadow_intermed_1 <= V_X_ANNUL_ALL_shadow;
		RIN_E_CTRL_ANNUL_intermed_1 <= RIN.E.CTRL.ANNUL;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_X_ANNUL_ALL_intermed_2 <= RIN_X_ANNUL_ALL_intermed_1;
		V_A_CTRL_ANNUL_shadow_intermed_1 <= V_A_CTRL_ANNUL_shadow;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_A_CTRL_ANNUL_intermed_2 <= RIN_A_CTRL_ANNUL_intermed_1;
		R_A_CTRL_ANNUL_intermed_1 <= R.A.CTRL.ANNUL;
		R_X_ANNUL_ALL_intermed_1 <= R.X.ANNUL_ALL;
		V_A_CTRL_RETT_shadow_intermed_1 <= V_A_CTRL_RETT_shadow;
		RIN_A_CTRL_RETT_intermed_1 <= RIN.A.CTRL.RETT;
		V_X_ANNUL_ALL_shadow_intermed_1 <= V_X_ANNUL_ALL_shadow;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_X_ANNUL_ALL_intermed_2 <= RIN_X_ANNUL_ALL_intermed_1;
		RIN_E_CTRL_RETT_intermed_1 <= RIN.E.CTRL.RETT;
		V_A_CTRL_ANNUL_shadow_intermed_1 <= V_A_CTRL_ANNUL_shadow;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_A_CTRL_ANNUL_intermed_2 <= RIN_A_CTRL_ANNUL_intermed_1;
		R_A_CTRL_ANNUL_intermed_1 <= R.A.CTRL.ANNUL;
		R_X_ANNUL_ALL_intermed_1 <= R.X.ANNUL_ALL;
		RIN_A_CTRL_WREG_intermed_1 <= RIN.A.CTRL.WREG;
		V_A_CTRL_WREG_shadow_intermed_1 <= V_A_CTRL_WREG_shadow;
		V_X_ANNUL_ALL_shadow_intermed_1 <= V_X_ANNUL_ALL_shadow;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_X_ANNUL_ALL_intermed_2 <= RIN_X_ANNUL_ALL_intermed_1;
		V_A_CTRL_ANNUL_shadow_intermed_1 <= V_A_CTRL_ANNUL_shadow;
		RIN_E_CTRL_WREG_intermed_1 <= RIN.E.CTRL.WREG;
		RIN_A_SU_intermed_1 <= RIN.A.SU;
		V_A_SU_shadow_intermed_1 <= V_A_SU_shadow;
		RIN_E_SU_intermed_1 <= RIN.E.SU;
		RIN_E_ET_intermed_1 <= RIN.E.ET;
		RIN_A_ET_intermed_1 <= RIN.A.ET;
		V_A_ET_shadow_intermed_1 <= V_A_ET_shadow;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_A_CTRL_ANNUL_intermed_2 <= RIN_A_CTRL_ANNUL_intermed_1;
		V_A_CTRL_WICC_shadow_intermed_1 <= V_A_CTRL_WICC_shadow;
		R_A_CTRL_ANNUL_intermed_1 <= R.A.CTRL.ANNUL;
		RIN_E_CTRL_WICC_intermed_1 <= RIN.E.CTRL.WICC;
		R_X_ANNUL_ALL_intermed_1 <= R.X.ANNUL_ALL;
		V_X_ANNUL_ALL_shadow_intermed_1 <= V_X_ANNUL_ALL_shadow;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_X_ANNUL_ALL_intermed_2 <= RIN_X_ANNUL_ALL_intermed_1;
		RIN_A_CTRL_WICC_intermed_1 <= RIN.A.CTRL.WICC;
		V_A_CTRL_ANNUL_shadow_intermed_1 <= V_A_CTRL_ANNUL_shadow;
		RIN_D_CWP_intermed_1 <= RIN.D.CWP;
		RIN_A_CWP_intermed_1 <= RIN.A.CWP;
		V_D_CWP_shadow_intermed_1 <= V_D_CWP_shadow;
		RIN_A_RFA1_intermed_1 <= RIN.A.RFA1;
		V_A_RFA1_shadow_intermed_1 <= V_A_RFA1_shadow;
		DBGI_DADDR9DOWNTO2_intermed_1 <= DBGI.DADDR ( 9 DOWNTO 2 );
		RIN_A_RFA1_intermed_1 <= RIN.A.RFA1;
		RIN_A_RFA2_intermed_1 <= RIN.A.RFA2;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_A_CTRL_WICC_intermed_1 <= RIN.A.CTRL.WICC;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_A_CTRL_WREG_intermed_1 <= RIN.A.CTRL.WREG;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_A_CTRL_RETT_intermed_1 <= RIN.A.CTRL.RETT;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_A_CTRL_WY_intermed_1 <= RIN.A.CTRL.WY;
		ICO_MEXC_intermed_1 <= ICO.MEXC;
		RIN_A_CTRL_TRAP_intermed_1 <= RIN.A.CTRL.TRAP;
		V_D_MEXC_shadow_intermed_1 <= V_D_MEXC_shadow;
		RIN_D_MEXC_intermed_1 <= RIN.D.MEXC;
		RIN_A_CTRL_TT_intermed_1 <= RIN.A.CTRL.TT;
		RIN_A_CTRL_INST_intermed_1 <= RIN.A.CTRL.INST;
		RIN_D_PC_intermed_1 <= RIN.D.PC;
		RIN_A_CTRL_PC_intermed_1 <= RIN.A.CTRL.PC;
		V_D_PC_shadow_intermed_1 <= V_D_PC_shadow;
		RIN_D_CNT_intermed_1 <= RIN.D.CNT;
		V_D_CNT_shadow_intermed_1 <= V_D_CNT_shadow;
		RIN_A_CTRL_CNT_intermed_1 <= RIN.A.CTRL.CNT;
		R_D_ANNUL_intermed_1 <= R.D.ANNUL;
		RIN_D_STEP_intermed_1 <= RIN.D.STEP;
		V_D_ANNUL_shadow_intermed_1 <= V_D_ANNUL_shadow;
		V_D_ANNUL_shadow_intermed_2 <= V_D_ANNUL_shadow_intermed_1;
		DBGI_STEP_intermed_1 <= DBGI.STEP;
		V_D_STEP_shadow_intermed_1 <= V_D_STEP_shadow;
		RIN_D_ANNUL_intermed_1 <= RIN.D.ANNUL;
		RIN_D_ANNUL_intermed_2 <= RIN_D_ANNUL_intermed_1;
		RIN_A_STEP_intermed_1 <= RIN.A.STEP;
		RIN_D_STEP_intermed_1 <= RIN.D.STEP;
		V_D_ANNUL_shadow_intermed_1 <= V_D_ANNUL_shadow;
		RIN_D_ANNUL_intermed_1 <= RIN.D.ANNUL;
		RIN_D_CNT_intermed_1 <= RIN.D.CNT;
		EX_ADD_RES32DOWNTO3_shadow_intermed_1 <= EX_ADD_RES32DOWNTO3_shadow;
		RIN_F_PC_intermed_1 <= RIN.F.PC;
		EX_JUMP_ADDRESS_shadow_intermed_1 <= EX_JUMP_ADDRESS_shadow;
		RIN_F_BRANCH_intermed_1 <= RIN.F.BRANCH;
		R_M_CTRL_PC31DOWNTO12_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 12 );
		R_M_CTRL_PC31DOWNTO12_intermed_2 <= R_M_CTRL_PC31DOWNTO12_intermed_1;
		R_M_CTRL_PC31DOWNTO12_intermed_3 <= R_M_CTRL_PC31DOWNTO12_intermed_2;
		V_D_PC31DOWNTO12_shadow_intermed_1 <= V_D_PC31DOWNTO12_shadow;
		V_D_PC31DOWNTO12_shadow_intermed_2 <= V_D_PC31DOWNTO12_shadow_intermed_1;
		V_D_PC31DOWNTO12_shadow_intermed_3 <= V_D_PC31DOWNTO12_shadow_intermed_2;
		V_D_PC31DOWNTO12_shadow_intermed_4 <= V_D_PC31DOWNTO12_shadow_intermed_3;
		V_D_PC31DOWNTO12_shadow_intermed_5 <= V_D_PC31DOWNTO12_shadow_intermed_4;
		V_D_PC31DOWNTO12_shadow_intermed_6 <= V_D_PC31DOWNTO12_shadow_intermed_5;
		V_D_PC31DOWNTO12_shadow_intermed_7 <= V_D_PC31DOWNTO12_shadow_intermed_6;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO12_shadow;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_4;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_6 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_5;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO12_shadow;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_3;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_5 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_4;
		EX_ADD_RES32DOWNTO330DOWNTO11_shadow_intermed_1 <= EX_ADD_RES32DOWNTO330DOWNTO11_shadow;
		EX_ADD_RES32DOWNTO330DOWNTO11_shadow_intermed_2 <= EX_ADD_RES32DOWNTO330DOWNTO11_shadow_intermed_1;
		RIN_F_PC31DOWNTO12_intermed_1 <= RIN.F.PC( 31 DOWNTO 12 );
		RIN_F_PC31DOWNTO12_intermed_2 <= RIN_F_PC31DOWNTO12_intermed_1;
		R_A_CTRL_PC31DOWNTO12_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 12 );
		R_A_CTRL_PC31DOWNTO12_intermed_2 <= R_A_CTRL_PC31DOWNTO12_intermed_1;
		R_A_CTRL_PC31DOWNTO12_intermed_3 <= R_A_CTRL_PC31DOWNTO12_intermed_2;
		R_A_CTRL_PC31DOWNTO12_intermed_4 <= R_A_CTRL_PC31DOWNTO12_intermed_3;
		R_A_CTRL_PC31DOWNTO12_intermed_5 <= R_A_CTRL_PC31DOWNTO12_intermed_4;
		R_E_CTRL_PC31DOWNTO12_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 12 );
		R_E_CTRL_PC31DOWNTO12_intermed_2 <= R_E_CTRL_PC31DOWNTO12_intermed_1;
		R_E_CTRL_PC31DOWNTO12_intermed_3 <= R_E_CTRL_PC31DOWNTO12_intermed_2;
		R_E_CTRL_PC31DOWNTO12_intermed_4 <= R_E_CTRL_PC31DOWNTO12_intermed_3;
		EX_JUMP_ADDRESS31DOWNTO12_shadow_intermed_1 <= EX_JUMP_ADDRESS31DOWNTO12_shadow;
		EX_JUMP_ADDRESS31DOWNTO12_shadow_intermed_2 <= EX_JUMP_ADDRESS31DOWNTO12_shadow_intermed_1;
		RIN_F_PC31DOWNTO12_intermed_1 <= RIN.F.PC ( 31 DOWNTO 12 );
		RIN_A_CTRL_PC31DOWNTO12_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 12 );
		RIN_A_CTRL_PC31DOWNTO12_intermed_2 <= RIN_A_CTRL_PC31DOWNTO12_intermed_1;
		RIN_A_CTRL_PC31DOWNTO12_intermed_3 <= RIN_A_CTRL_PC31DOWNTO12_intermed_2;
		RIN_A_CTRL_PC31DOWNTO12_intermed_4 <= RIN_A_CTRL_PC31DOWNTO12_intermed_3;
		RIN_A_CTRL_PC31DOWNTO12_intermed_5 <= RIN_A_CTRL_PC31DOWNTO12_intermed_4;
		RIN_A_CTRL_PC31DOWNTO12_intermed_6 <= RIN_A_CTRL_PC31DOWNTO12_intermed_5;
		RIN_E_CTRL_PC31DOWNTO12_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 12 );
		RIN_E_CTRL_PC31DOWNTO12_intermed_2 <= RIN_E_CTRL_PC31DOWNTO12_intermed_1;
		RIN_E_CTRL_PC31DOWNTO12_intermed_3 <= RIN_E_CTRL_PC31DOWNTO12_intermed_2;
		RIN_E_CTRL_PC31DOWNTO12_intermed_4 <= RIN_E_CTRL_PC31DOWNTO12_intermed_3;
		RIN_E_CTRL_PC31DOWNTO12_intermed_5 <= RIN_E_CTRL_PC31DOWNTO12_intermed_4;
		V_F_PC31DOWNTO12_shadow_intermed_1 <= V_F_PC31DOWNTO12_shadow;
		V_F_PC31DOWNTO12_shadow_intermed_2 <= V_F_PC31DOWNTO12_shadow_intermed_1;
		IRIN_ADDR31DOWNTO12_intermed_1 <= IRIN.ADDR( 31 DOWNTO 12 );
		IRIN_ADDR31DOWNTO12_intermed_2 <= IRIN_ADDR31DOWNTO12_intermed_1;
		V_X_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO12_shadow;
		V_X_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_X_CTRL_PC31DOWNTO12_shadow_intermed_2;
		EX_ADD_RES32DOWNTO332DOWNTO13_shadow_intermed_1 <= EX_ADD_RES32DOWNTO332DOWNTO13_shadow;
		EX_ADD_RES32DOWNTO332DOWNTO13_shadow_intermed_2 <= EX_ADD_RES32DOWNTO332DOWNTO13_shadow_intermed_1;
		XC_TRAP_ADDRESS31DOWNTO12_shadow_intermed_1 <= XC_TRAP_ADDRESS31DOWNTO12_shadow;
		R_F_PC31DOWNTO12_intermed_1 <= R.F.PC( 31 DOWNTO 12 );
		RIN_M_CTRL_PC31DOWNTO12_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 12 );
		RIN_M_CTRL_PC31DOWNTO12_intermed_2 <= RIN_M_CTRL_PC31DOWNTO12_intermed_1;
		RIN_M_CTRL_PC31DOWNTO12_intermed_3 <= RIN_M_CTRL_PC31DOWNTO12_intermed_2;
		RIN_M_CTRL_PC31DOWNTO12_intermed_4 <= RIN_M_CTRL_PC31DOWNTO12_intermed_3;
		IR_ADDR31DOWNTO12_intermed_1 <= IR.ADDR( 31 DOWNTO 12 );
		R_X_CTRL_PC31DOWNTO12_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 12 );
		R_X_CTRL_PC31DOWNTO12_intermed_2 <= R_X_CTRL_PC31DOWNTO12_intermed_1;
		R_D_PC31DOWNTO12_intermed_1 <= R.D.PC( 31 DOWNTO 12 );
		R_D_PC31DOWNTO12_intermed_2 <= R_D_PC31DOWNTO12_intermed_1;
		R_D_PC31DOWNTO12_intermed_3 <= R_D_PC31DOWNTO12_intermed_2;
		R_D_PC31DOWNTO12_intermed_4 <= R_D_PC31DOWNTO12_intermed_3;
		R_D_PC31DOWNTO12_intermed_5 <= R_D_PC31DOWNTO12_intermed_4;
		R_D_PC31DOWNTO12_intermed_6 <= R_D_PC31DOWNTO12_intermed_5;
		RIN_X_CTRL_PC31DOWNTO12_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 12 );
		RIN_X_CTRL_PC31DOWNTO12_intermed_2 <= RIN_X_CTRL_PC31DOWNTO12_intermed_1;
		RIN_X_CTRL_PC31DOWNTO12_intermed_3 <= RIN_X_CTRL_PC31DOWNTO12_intermed_2;
		RIN_D_PC31DOWNTO12_intermed_1 <= RIN.D.PC( 31 DOWNTO 12 );
		RIN_D_PC31DOWNTO12_intermed_2 <= RIN_D_PC31DOWNTO12_intermed_1;
		RIN_D_PC31DOWNTO12_intermed_3 <= RIN_D_PC31DOWNTO12_intermed_2;
		RIN_D_PC31DOWNTO12_intermed_4 <= RIN_D_PC31DOWNTO12_intermed_3;
		RIN_D_PC31DOWNTO12_intermed_5 <= RIN_D_PC31DOWNTO12_intermed_4;
		RIN_D_PC31DOWNTO12_intermed_6 <= RIN_D_PC31DOWNTO12_intermed_5;
		RIN_D_PC31DOWNTO12_intermed_7 <= RIN_D_PC31DOWNTO12_intermed_6;
		VIR_ADDR31DOWNTO12_shadow_intermed_1 <= VIR_ADDR31DOWNTO12_shadow;
		VIR_ADDR31DOWNTO12_shadow_intermed_2 <= VIR_ADDR31DOWNTO12_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO12_shadow;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_4 <= V_M_CTRL_PC31DOWNTO12_shadow_intermed_3;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_3 <= RIN_M_CTRL_PC31DOWNTO2_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_4 <= RIN_M_CTRL_PC31DOWNTO2_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_5 <= V_D_PC31DOWNTO2_shadow_intermed_4;
		V_D_PC31DOWNTO2_shadow_intermed_6 <= V_D_PC31DOWNTO2_shadow_intermed_5;
		V_D_PC31DOWNTO2_shadow_intermed_7 <= V_D_PC31DOWNTO2_shadow_intermed_6;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_5 <= RIN_D_PC31DOWNTO2_intermed_4;
		RIN_D_PC31DOWNTO2_intermed_6 <= RIN_D_PC31DOWNTO2_intermed_5;
		RIN_D_PC31DOWNTO2_intermed_7 <= RIN_D_PC31DOWNTO2_intermed_6;
		EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_1 <= EX_ADD_RES32DOWNTO332DOWNTO3_shadow;
		EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_2 <= EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_1;
		V_F_PC31DOWNTO2_shadow_intermed_1 <= V_F_PC31DOWNTO2_shadow;
		V_F_PC31DOWNTO2_shadow_intermed_2 <= V_F_PC31DOWNTO2_shadow_intermed_1;
		RIN_F_PC31DOWNTO2_intermed_1 <= RIN.F.PC( 31 DOWNTO 2 );
		RIN_F_PC31DOWNTO2_intermed_2 <= RIN_F_PC31DOWNTO2_intermed_1;
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_2 <= RIN_X_CTRL_PC31DOWNTO2_intermed_1;
		RIN_X_CTRL_PC31DOWNTO2_intermed_3 <= RIN_X_CTRL_PC31DOWNTO2_intermed_2;
		IRIN_ADDR31DOWNTO2_intermed_1 <= IRIN.ADDR( 31 DOWNTO 2 );
		IRIN_ADDR31DOWNTO2_intermed_2 <= IRIN_ADDR31DOWNTO2_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_6 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_5;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		R_D_PC31DOWNTO2_intermed_4 <= R_D_PC31DOWNTO2_intermed_3;
		R_D_PC31DOWNTO2_intermed_5 <= R_D_PC31DOWNTO2_intermed_4;
		R_D_PC31DOWNTO2_intermed_6 <= R_D_PC31DOWNTO2_intermed_5;
		R_F_PC31DOWNTO2_intermed_1 <= R.F.PC( 31 DOWNTO 2 );
		VIR_ADDR31DOWNTO2_shadow_intermed_1 <= VIR_ADDR31DOWNTO2_shadow;
		VIR_ADDR31DOWNTO2_shadow_intermed_2 <= VIR_ADDR31DOWNTO2_shadow_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 2 );
		R_M_CTRL_PC31DOWNTO2_intermed_2 <= R_M_CTRL_PC31DOWNTO2_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_3 <= R_M_CTRL_PC31DOWNTO2_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_4;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		RIN_A_CTRL_PC31DOWNTO2_intermed_5 <= RIN_A_CTRL_PC31DOWNTO2_intermed_4;
		RIN_A_CTRL_PC31DOWNTO2_intermed_6 <= RIN_A_CTRL_PC31DOWNTO2_intermed_5;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_4 <= R_A_CTRL_PC31DOWNTO2_intermed_3;
		R_A_CTRL_PC31DOWNTO2_intermed_5 <= R_A_CTRL_PC31DOWNTO2_intermed_4;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_3;
		R_X_CTRL_PC31DOWNTO2_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 2 );
		R_X_CTRL_PC31DOWNTO2_intermed_2 <= R_X_CTRL_PC31DOWNTO2_intermed_1;
		XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_1 <= XC_TRAP_ADDRESS31DOWNTO2_shadow;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_3 <= R_E_CTRL_PC31DOWNTO2_intermed_2;
		R_E_CTRL_PC31DOWNTO2_intermed_4 <= R_E_CTRL_PC31DOWNTO2_intermed_3;
		EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_1 <= EX_JUMP_ADDRESS31DOWNTO2_shadow;
		EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_2 <= EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_1;
		RIN_F_PC31DOWNTO2_intermed_1 <= RIN.F.PC ( 31 DOWNTO 2 );
		IR_ADDR31DOWNTO2_intermed_1 <= IR.ADDR( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_4 <= RIN_E_CTRL_PC31DOWNTO2_intermed_3;
		RIN_E_CTRL_PC31DOWNTO2_intermed_5 <= RIN_E_CTRL_PC31DOWNTO2_intermed_4;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO2_shadow;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_3 <= RIN_M_CTRL_PC31DOWNTO2_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_4 <= RIN_M_CTRL_PC31DOWNTO2_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_5 <= V_D_PC31DOWNTO2_shadow_intermed_4;
		V_D_PC31DOWNTO2_shadow_intermed_6 <= V_D_PC31DOWNTO2_shadow_intermed_5;
		V_D_PC31DOWNTO2_shadow_intermed_7 <= V_D_PC31DOWNTO2_shadow_intermed_6;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_5 <= RIN_D_PC31DOWNTO2_intermed_4;
		RIN_D_PC31DOWNTO2_intermed_6 <= RIN_D_PC31DOWNTO2_intermed_5;
		RIN_D_PC31DOWNTO2_intermed_7 <= RIN_D_PC31DOWNTO2_intermed_6;
		EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_1 <= EX_ADD_RES32DOWNTO332DOWNTO3_shadow;
		V_F_PC31DOWNTO2_shadow_intermed_1 <= V_F_PC31DOWNTO2_shadow;
		RIN_F_PC31DOWNTO2_intermed_1 <= RIN.F.PC( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_2 <= RIN_X_CTRL_PC31DOWNTO2_intermed_1;
		RIN_X_CTRL_PC31DOWNTO2_intermed_3 <= RIN_X_CTRL_PC31DOWNTO2_intermed_2;
		IRIN_ADDR31DOWNTO2_intermed_1 <= IRIN.ADDR( 31 DOWNTO 2 );
		IRIN_ADDR31DOWNTO2_intermed_2 <= IRIN_ADDR31DOWNTO2_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_6 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_5;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		R_D_PC31DOWNTO2_intermed_4 <= R_D_PC31DOWNTO2_intermed_3;
		R_D_PC31DOWNTO2_intermed_5 <= R_D_PC31DOWNTO2_intermed_4;
		R_D_PC31DOWNTO2_intermed_6 <= R_D_PC31DOWNTO2_intermed_5;
		VIR_ADDR31DOWNTO2_shadow_intermed_1 <= VIR_ADDR31DOWNTO2_shadow;
		VIR_ADDR31DOWNTO2_shadow_intermed_2 <= VIR_ADDR31DOWNTO2_shadow_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 2 );
		R_M_CTRL_PC31DOWNTO2_intermed_2 <= R_M_CTRL_PC31DOWNTO2_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_3 <= R_M_CTRL_PC31DOWNTO2_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_4;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		RIN_A_CTRL_PC31DOWNTO2_intermed_5 <= RIN_A_CTRL_PC31DOWNTO2_intermed_4;
		RIN_A_CTRL_PC31DOWNTO2_intermed_6 <= RIN_A_CTRL_PC31DOWNTO2_intermed_5;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_4 <= R_A_CTRL_PC31DOWNTO2_intermed_3;
		R_A_CTRL_PC31DOWNTO2_intermed_5 <= R_A_CTRL_PC31DOWNTO2_intermed_4;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_3;
		R_X_CTRL_PC31DOWNTO2_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 2 );
		R_X_CTRL_PC31DOWNTO2_intermed_2 <= R_X_CTRL_PC31DOWNTO2_intermed_1;
		XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_1 <= XC_TRAP_ADDRESS31DOWNTO2_shadow;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_3 <= R_E_CTRL_PC31DOWNTO2_intermed_2;
		R_E_CTRL_PC31DOWNTO2_intermed_4 <= R_E_CTRL_PC31DOWNTO2_intermed_3;
		EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_1 <= EX_JUMP_ADDRESS31DOWNTO2_shadow;
		IR_ADDR31DOWNTO2_intermed_1 <= IR.ADDR( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_4 <= RIN_E_CTRL_PC31DOWNTO2_intermed_3;
		RIN_E_CTRL_PC31DOWNTO2_intermed_5 <= RIN_E_CTRL_PC31DOWNTO2_intermed_4;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO2_shadow;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_2;
		RIN_D_INST0_intermed_1 <= RIN.D.INST ( 0 );
		R_D_INST0_intermed_1 <= R.D.INST( 0 );
		V_D_INST0_shadow_intermed_1 <= V_D_INST0_shadow;
		V_D_INST0_shadow_intermed_2 <= V_D_INST0_shadow_intermed_1;
		RIN_D_INST0_intermed_1 <= RIN.D.INST( 0 );
		RIN_D_INST0_intermed_2 <= RIN_D_INST0_intermed_1;
		RIN_D_INST1_intermed_1 <= RIN.D.INST ( 1 );
		R_D_INST1_intermed_1 <= R.D.INST( 1 );
		V_D_INST1_shadow_intermed_1 <= V_D_INST1_shadow;
		V_D_INST1_shadow_intermed_2 <= V_D_INST1_shadow_intermed_1;
		RIN_D_INST1_intermed_1 <= RIN.D.INST( 1 );
		RIN_D_INST1_intermed_2 <= RIN_D_INST1_intermed_1;
		RIN_D_SET_intermed_1 <= RIN.D.SET;
		RIN_D_MEXC_intermed_1 <= RIN.D.MEXC;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA ( 0 )( 31 );
		RIN_E_OP131_intermed_1 <= RIN.E.OP1( 31 );
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_2 <= V_X_DATA031_shadow_intermed_1;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA( 0 )( 31 );
		RIN_X_DATA031_intermed_2 <= RIN_X_DATA031_intermed_1;
		DCO_DATA031_intermed_1 <= DCO.DATA ( 0 )( 31 );
		V_E_OP131_shadow_intermed_1 <= V_E_OP131_shadow;
		R_X_DATA031_intermed_1 <= R.X.DATA( 0 )( 31 );
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA ( 0 )( 31 );
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_2 <= V_X_DATA031_shadow_intermed_1;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA( 0 )( 31 );
		RIN_X_DATA031_intermed_2 <= RIN_X_DATA031_intermed_1;
		DCO_DATA031_intermed_1 <= DCO.DATA ( 0 )( 31 );
		RIN_E_OP231_intermed_1 <= RIN.E.OP2( 31 );
		R_X_DATA031_intermed_1 <= R.X.DATA( 0 )( 31 );
		V_E_OP231_shadow_intermed_1 <= V_E_OP231_shadow;
		V_D_ANNUL_shadow_intermed_1 <= V_D_ANNUL_shadow;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_D_ANNUL_intermed_1 <= RIN.D.ANNUL;
		V_X_DATA03_shadow_intermed_1 <= V_X_DATA03_shadow;
		V_X_DATA03_shadow_intermed_2 <= V_X_DATA03_shadow_intermed_1;
		V_X_DATA03_shadow_intermed_1 <= V_X_DATA03_shadow;
		DCO_DATA03_intermed_1 <= DCO.DATA ( 0 )( 3 );
		RIN_X_DATA03_intermed_1 <= RIN.X.DATA ( 0 )( 3 );
		R_X_DATA03_intermed_1 <= R.X.DATA( 0 )( 3 );
		RIN_X_DATA03_intermed_1 <= RIN.X.DATA( 0 )( 3 );
		RIN_X_DATA03_intermed_2 <= RIN_X_DATA03_intermed_1;
		RIN_E_OP13_intermed_1 <= RIN.E.OP1( 3 );
		V_E_OP13_shadow_intermed_1 <= V_E_OP13_shadow;
		V_X_DATA03_shadow_intermed_1 <= V_X_DATA03_shadow;
		V_X_DATA03_shadow_intermed_2 <= V_X_DATA03_shadow_intermed_1;
		V_X_DATA03_shadow_intermed_1 <= V_X_DATA03_shadow;
		DCO_DATA03_intermed_1 <= DCO.DATA ( 0 )( 3 );
		RIN_X_DATA03_intermed_1 <= RIN.X.DATA ( 0 )( 3 );
		R_X_DATA03_intermed_1 <= R.X.DATA( 0 )( 3 );
		RIN_X_DATA03_intermed_1 <= RIN.X.DATA( 0 )( 3 );
		RIN_X_DATA03_intermed_2 <= RIN_X_DATA03_intermed_1;
		RIN_E_OP23_intermed_1 <= RIN.E.OP2( 3 );
		V_E_OP23_shadow_intermed_1 <= V_E_OP23_shadow;
		R_M_CTRL_PC31DOWNTO12_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 12 );
		R_M_CTRL_PC31DOWNTO12_intermed_2 <= R_M_CTRL_PC31DOWNTO12_intermed_1;
		R_M_CTRL_PC31DOWNTO12_intermed_3 <= R_M_CTRL_PC31DOWNTO12_intermed_2;
		V_D_PC31DOWNTO12_shadow_intermed_1 <= V_D_PC31DOWNTO12_shadow;
		V_D_PC31DOWNTO12_shadow_intermed_2 <= V_D_PC31DOWNTO12_shadow_intermed_1;
		V_D_PC31DOWNTO12_shadow_intermed_3 <= V_D_PC31DOWNTO12_shadow_intermed_2;
		V_D_PC31DOWNTO12_shadow_intermed_4 <= V_D_PC31DOWNTO12_shadow_intermed_3;
		V_D_PC31DOWNTO12_shadow_intermed_5 <= V_D_PC31DOWNTO12_shadow_intermed_4;
		V_D_PC31DOWNTO12_shadow_intermed_6 <= V_D_PC31DOWNTO12_shadow_intermed_5;
		V_D_PC31DOWNTO12_shadow_intermed_7 <= V_D_PC31DOWNTO12_shadow_intermed_6;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO12_shadow;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_4;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_6 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_5;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO12_shadow;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_3;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_5 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_4;
		EX_ADD_RES32DOWNTO330DOWNTO11_shadow_intermed_1 <= EX_ADD_RES32DOWNTO330DOWNTO11_shadow;
		RIN_F_PC31DOWNTO12_intermed_1 <= RIN.F.PC( 31 DOWNTO 12 );
		R_A_CTRL_PC31DOWNTO12_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 12 );
		R_A_CTRL_PC31DOWNTO12_intermed_2 <= R_A_CTRL_PC31DOWNTO12_intermed_1;
		R_A_CTRL_PC31DOWNTO12_intermed_3 <= R_A_CTRL_PC31DOWNTO12_intermed_2;
		R_A_CTRL_PC31DOWNTO12_intermed_4 <= R_A_CTRL_PC31DOWNTO12_intermed_3;
		R_A_CTRL_PC31DOWNTO12_intermed_5 <= R_A_CTRL_PC31DOWNTO12_intermed_4;
		R_E_CTRL_PC31DOWNTO12_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 12 );
		R_E_CTRL_PC31DOWNTO12_intermed_2 <= R_E_CTRL_PC31DOWNTO12_intermed_1;
		R_E_CTRL_PC31DOWNTO12_intermed_3 <= R_E_CTRL_PC31DOWNTO12_intermed_2;
		R_E_CTRL_PC31DOWNTO12_intermed_4 <= R_E_CTRL_PC31DOWNTO12_intermed_3;
		EX_JUMP_ADDRESS31DOWNTO12_shadow_intermed_1 <= EX_JUMP_ADDRESS31DOWNTO12_shadow;
		RIN_A_CTRL_PC31DOWNTO12_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 12 );
		RIN_A_CTRL_PC31DOWNTO12_intermed_2 <= RIN_A_CTRL_PC31DOWNTO12_intermed_1;
		RIN_A_CTRL_PC31DOWNTO12_intermed_3 <= RIN_A_CTRL_PC31DOWNTO12_intermed_2;
		RIN_A_CTRL_PC31DOWNTO12_intermed_4 <= RIN_A_CTRL_PC31DOWNTO12_intermed_3;
		RIN_A_CTRL_PC31DOWNTO12_intermed_5 <= RIN_A_CTRL_PC31DOWNTO12_intermed_4;
		RIN_A_CTRL_PC31DOWNTO12_intermed_6 <= RIN_A_CTRL_PC31DOWNTO12_intermed_5;
		RIN_E_CTRL_PC31DOWNTO12_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 12 );
		RIN_E_CTRL_PC31DOWNTO12_intermed_2 <= RIN_E_CTRL_PC31DOWNTO12_intermed_1;
		RIN_E_CTRL_PC31DOWNTO12_intermed_3 <= RIN_E_CTRL_PC31DOWNTO12_intermed_2;
		RIN_E_CTRL_PC31DOWNTO12_intermed_4 <= RIN_E_CTRL_PC31DOWNTO12_intermed_3;
		RIN_E_CTRL_PC31DOWNTO12_intermed_5 <= RIN_E_CTRL_PC31DOWNTO12_intermed_4;
		V_F_PC31DOWNTO12_shadow_intermed_1 <= V_F_PC31DOWNTO12_shadow;
		IRIN_ADDR31DOWNTO12_intermed_1 <= IRIN.ADDR( 31 DOWNTO 12 );
		IRIN_ADDR31DOWNTO12_intermed_2 <= IRIN_ADDR31DOWNTO12_intermed_1;
		V_X_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO12_shadow;
		V_X_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_X_CTRL_PC31DOWNTO12_shadow_intermed_2;
		EX_ADD_RES32DOWNTO332DOWNTO13_shadow_intermed_1 <= EX_ADD_RES32DOWNTO332DOWNTO13_shadow;
		RIN_M_CTRL_PC31DOWNTO12_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 12 );
		RIN_M_CTRL_PC31DOWNTO12_intermed_2 <= RIN_M_CTRL_PC31DOWNTO12_intermed_1;
		RIN_M_CTRL_PC31DOWNTO12_intermed_3 <= RIN_M_CTRL_PC31DOWNTO12_intermed_2;
		RIN_M_CTRL_PC31DOWNTO12_intermed_4 <= RIN_M_CTRL_PC31DOWNTO12_intermed_3;
		IR_ADDR31DOWNTO12_intermed_1 <= IR.ADDR( 31 DOWNTO 12 );
		R_X_CTRL_PC31DOWNTO12_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 12 );
		R_X_CTRL_PC31DOWNTO12_intermed_2 <= R_X_CTRL_PC31DOWNTO12_intermed_1;
		R_D_PC31DOWNTO12_intermed_1 <= R.D.PC( 31 DOWNTO 12 );
		R_D_PC31DOWNTO12_intermed_2 <= R_D_PC31DOWNTO12_intermed_1;
		R_D_PC31DOWNTO12_intermed_3 <= R_D_PC31DOWNTO12_intermed_2;
		R_D_PC31DOWNTO12_intermed_4 <= R_D_PC31DOWNTO12_intermed_3;
		R_D_PC31DOWNTO12_intermed_5 <= R_D_PC31DOWNTO12_intermed_4;
		R_D_PC31DOWNTO12_intermed_6 <= R_D_PC31DOWNTO12_intermed_5;
		RIN_X_CTRL_PC31DOWNTO12_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 12 );
		RIN_X_CTRL_PC31DOWNTO12_intermed_2 <= RIN_X_CTRL_PC31DOWNTO12_intermed_1;
		RIN_X_CTRL_PC31DOWNTO12_intermed_3 <= RIN_X_CTRL_PC31DOWNTO12_intermed_2;
		RIN_D_PC31DOWNTO12_intermed_1 <= RIN.D.PC( 31 DOWNTO 12 );
		RIN_D_PC31DOWNTO12_intermed_2 <= RIN_D_PC31DOWNTO12_intermed_1;
		RIN_D_PC31DOWNTO12_intermed_3 <= RIN_D_PC31DOWNTO12_intermed_2;
		RIN_D_PC31DOWNTO12_intermed_4 <= RIN_D_PC31DOWNTO12_intermed_3;
		RIN_D_PC31DOWNTO12_intermed_5 <= RIN_D_PC31DOWNTO12_intermed_4;
		RIN_D_PC31DOWNTO12_intermed_6 <= RIN_D_PC31DOWNTO12_intermed_5;
		RIN_D_PC31DOWNTO12_intermed_7 <= RIN_D_PC31DOWNTO12_intermed_6;
		VIR_ADDR31DOWNTO12_shadow_intermed_1 <= VIR_ADDR31DOWNTO12_shadow;
		VIR_ADDR31DOWNTO12_shadow_intermed_2 <= VIR_ADDR31DOWNTO12_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO12_shadow;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_4 <= V_M_CTRL_PC31DOWNTO12_shadow_intermed_3;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_3 <= RIN_M_CTRL_PC31DOWNTO2_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_4 <= RIN_M_CTRL_PC31DOWNTO2_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_5 <= V_D_PC31DOWNTO2_shadow_intermed_4;
		V_D_PC31DOWNTO2_shadow_intermed_6 <= V_D_PC31DOWNTO2_shadow_intermed_5;
		V_D_PC31DOWNTO2_shadow_intermed_7 <= V_D_PC31DOWNTO2_shadow_intermed_6;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_5 <= RIN_D_PC31DOWNTO2_intermed_4;
		RIN_D_PC31DOWNTO2_intermed_6 <= RIN_D_PC31DOWNTO2_intermed_5;
		RIN_D_PC31DOWNTO2_intermed_7 <= RIN_D_PC31DOWNTO2_intermed_6;
		EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_1 <= EX_ADD_RES32DOWNTO332DOWNTO3_shadow;
		V_F_PC31DOWNTO2_shadow_intermed_1 <= V_F_PC31DOWNTO2_shadow;
		RIN_F_PC31DOWNTO2_intermed_1 <= RIN.F.PC( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_2 <= RIN_X_CTRL_PC31DOWNTO2_intermed_1;
		RIN_X_CTRL_PC31DOWNTO2_intermed_3 <= RIN_X_CTRL_PC31DOWNTO2_intermed_2;
		IRIN_ADDR31DOWNTO2_intermed_1 <= IRIN.ADDR( 31 DOWNTO 2 );
		IRIN_ADDR31DOWNTO2_intermed_2 <= IRIN_ADDR31DOWNTO2_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_6 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_5;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		R_D_PC31DOWNTO2_intermed_4 <= R_D_PC31DOWNTO2_intermed_3;
		R_D_PC31DOWNTO2_intermed_5 <= R_D_PC31DOWNTO2_intermed_4;
		R_D_PC31DOWNTO2_intermed_6 <= R_D_PC31DOWNTO2_intermed_5;
		VIR_ADDR31DOWNTO2_shadow_intermed_1 <= VIR_ADDR31DOWNTO2_shadow;
		VIR_ADDR31DOWNTO2_shadow_intermed_2 <= VIR_ADDR31DOWNTO2_shadow_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 2 );
		R_M_CTRL_PC31DOWNTO2_intermed_2 <= R_M_CTRL_PC31DOWNTO2_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_3 <= R_M_CTRL_PC31DOWNTO2_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_4;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		RIN_A_CTRL_PC31DOWNTO2_intermed_5 <= RIN_A_CTRL_PC31DOWNTO2_intermed_4;
		RIN_A_CTRL_PC31DOWNTO2_intermed_6 <= RIN_A_CTRL_PC31DOWNTO2_intermed_5;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_4 <= R_A_CTRL_PC31DOWNTO2_intermed_3;
		R_A_CTRL_PC31DOWNTO2_intermed_5 <= R_A_CTRL_PC31DOWNTO2_intermed_4;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_3;
		R_X_CTRL_PC31DOWNTO2_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 2 );
		R_X_CTRL_PC31DOWNTO2_intermed_2 <= R_X_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_3 <= R_E_CTRL_PC31DOWNTO2_intermed_2;
		R_E_CTRL_PC31DOWNTO2_intermed_4 <= R_E_CTRL_PC31DOWNTO2_intermed_3;
		EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_1 <= EX_JUMP_ADDRESS31DOWNTO2_shadow;
		IR_ADDR31DOWNTO2_intermed_1 <= IR.ADDR( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_4 <= RIN_E_CTRL_PC31DOWNTO2_intermed_3;
		RIN_E_CTRL_PC31DOWNTO2_intermed_5 <= RIN_E_CTRL_PC31DOWNTO2_intermed_4;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO2_shadow;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_3 <= RIN_M_CTRL_PC31DOWNTO2_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_4 <= RIN_M_CTRL_PC31DOWNTO2_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_5 <= V_D_PC31DOWNTO2_shadow_intermed_4;
		V_D_PC31DOWNTO2_shadow_intermed_6 <= V_D_PC31DOWNTO2_shadow_intermed_5;
		V_D_PC31DOWNTO2_shadow_intermed_7 <= V_D_PC31DOWNTO2_shadow_intermed_6;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_5 <= RIN_D_PC31DOWNTO2_intermed_4;
		RIN_D_PC31DOWNTO2_intermed_6 <= RIN_D_PC31DOWNTO2_intermed_5;
		RIN_D_PC31DOWNTO2_intermed_7 <= RIN_D_PC31DOWNTO2_intermed_6;
		EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_1 <= EX_ADD_RES32DOWNTO332DOWNTO3_shadow;
		RIN_F_PC31DOWNTO2_intermed_1 <= RIN.F.PC( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_2 <= RIN_X_CTRL_PC31DOWNTO2_intermed_1;
		RIN_X_CTRL_PC31DOWNTO2_intermed_3 <= RIN_X_CTRL_PC31DOWNTO2_intermed_2;
		IRIN_ADDR31DOWNTO2_intermed_1 <= IRIN.ADDR( 31 DOWNTO 2 );
		IRIN_ADDR31DOWNTO2_intermed_2 <= IRIN_ADDR31DOWNTO2_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_6 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_5;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		R_D_PC31DOWNTO2_intermed_4 <= R_D_PC31DOWNTO2_intermed_3;
		R_D_PC31DOWNTO2_intermed_5 <= R_D_PC31DOWNTO2_intermed_4;
		R_D_PC31DOWNTO2_intermed_6 <= R_D_PC31DOWNTO2_intermed_5;
		VIR_ADDR31DOWNTO2_shadow_intermed_1 <= VIR_ADDR31DOWNTO2_shadow;
		VIR_ADDR31DOWNTO2_shadow_intermed_2 <= VIR_ADDR31DOWNTO2_shadow_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 2 );
		R_M_CTRL_PC31DOWNTO2_intermed_2 <= R_M_CTRL_PC31DOWNTO2_intermed_1;
		R_M_CTRL_PC31DOWNTO2_intermed_3 <= R_M_CTRL_PC31DOWNTO2_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_4;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		RIN_A_CTRL_PC31DOWNTO2_intermed_5 <= RIN_A_CTRL_PC31DOWNTO2_intermed_4;
		RIN_A_CTRL_PC31DOWNTO2_intermed_6 <= RIN_A_CTRL_PC31DOWNTO2_intermed_5;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_4 <= R_A_CTRL_PC31DOWNTO2_intermed_3;
		R_A_CTRL_PC31DOWNTO2_intermed_5 <= R_A_CTRL_PC31DOWNTO2_intermed_4;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_3;
		R_X_CTRL_PC31DOWNTO2_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 2 );
		R_X_CTRL_PC31DOWNTO2_intermed_2 <= R_X_CTRL_PC31DOWNTO2_intermed_1;
		XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_1 <= XC_TRAP_ADDRESS31DOWNTO2_shadow;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_3 <= R_E_CTRL_PC31DOWNTO2_intermed_2;
		R_E_CTRL_PC31DOWNTO2_intermed_4 <= R_E_CTRL_PC31DOWNTO2_intermed_3;
		EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_1 <= EX_JUMP_ADDRESS31DOWNTO2_shadow;
		IR_ADDR31DOWNTO2_intermed_1 <= IR.ADDR( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_4 <= RIN_E_CTRL_PC31DOWNTO2_intermed_3;
		RIN_E_CTRL_PC31DOWNTO2_intermed_5 <= RIN_E_CTRL_PC31DOWNTO2_intermed_4;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO2_shadow;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_2;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA ( 0 )( 31 );
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_2 <= V_X_DATA031_shadow_intermed_1;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA( 0 )( 31 );
		RIN_X_DATA031_intermed_2 <= RIN_X_DATA031_intermed_1;
		DCO_DATA031_intermed_1 <= DCO.DATA ( 0 )( 31 );
		RIN_E_OP231_intermed_1 <= RIN.E.OP2( 31 );
		R_X_DATA031_intermed_1 <= R.X.DATA( 0 )( 31 );
		V_E_OP231_shadow_intermed_1 <= V_E_OP231_shadow;
		V_M_CTRL_RD7DOWNTO0_shadow_intermed_1 <= V_M_CTRL_RD7DOWNTO0_shadow;
		V_M_CTRL_RD7DOWNTO0_shadow_intermed_2 <= V_M_CTRL_RD7DOWNTO0_shadow_intermed_1;
		V_E_CTRL_RD7DOWNTO0_shadow_intermed_1 <= V_E_CTRL_RD7DOWNTO0_shadow;
		V_E_CTRL_RD7DOWNTO0_shadow_intermed_2 <= V_E_CTRL_RD7DOWNTO0_shadow_intermed_1;
		V_E_CTRL_RD7DOWNTO0_shadow_intermed_3 <= V_E_CTRL_RD7DOWNTO0_shadow_intermed_2;
		R_E_CTRL_RD7DOWNTO0_intermed_1 <= R.E.CTRL.RD ( 7 DOWNTO 0 );
		R_E_CTRL_RD7DOWNTO0_intermed_2 <= R_E_CTRL_RD7DOWNTO0_intermed_1;
		V_A_CTRL_RD7DOWNTO0_shadow_intermed_1 <= V_A_CTRL_RD7DOWNTO0_shadow;
		V_A_CTRL_RD7DOWNTO0_shadow_intermed_2 <= V_A_CTRL_RD7DOWNTO0_shadow_intermed_1;
		V_A_CTRL_RD7DOWNTO0_shadow_intermed_3 <= V_A_CTRL_RD7DOWNTO0_shadow_intermed_2;
		V_A_CTRL_RD7DOWNTO0_shadow_intermed_4 <= V_A_CTRL_RD7DOWNTO0_shadow_intermed_3;
		RIN_A_CTRL_RD7DOWNTO0_intermed_1 <= RIN.A.CTRL.RD ( 7 DOWNTO 0 );
		RIN_A_CTRL_RD7DOWNTO0_intermed_2 <= RIN_A_CTRL_RD7DOWNTO0_intermed_1;
		RIN_A_CTRL_RD7DOWNTO0_intermed_3 <= RIN_A_CTRL_RD7DOWNTO0_intermed_2;
		RIN_A_CTRL_RD7DOWNTO0_intermed_4 <= RIN_A_CTRL_RD7DOWNTO0_intermed_3;
		R_M_CTRL_RD7DOWNTO0_intermed_1 <= R.M.CTRL.RD ( 7 DOWNTO 0 );
		R_A_CTRL_RD7DOWNTO0_intermed_1 <= R.A.CTRL.RD ( 7 DOWNTO 0 );
		R_A_CTRL_RD7DOWNTO0_intermed_2 <= R_A_CTRL_RD7DOWNTO0_intermed_1;
		R_A_CTRL_RD7DOWNTO0_intermed_3 <= R_A_CTRL_RD7DOWNTO0_intermed_2;
		RIN_E_CTRL_RD7DOWNTO0_intermed_1 <= RIN.E.CTRL.RD ( 7 DOWNTO 0 );
		RIN_E_CTRL_RD7DOWNTO0_intermed_2 <= RIN_E_CTRL_RD7DOWNTO0_intermed_1;
		RIN_E_CTRL_RD7DOWNTO0_intermed_3 <= RIN_E_CTRL_RD7DOWNTO0_intermed_2;
		RIN_X_CTRL_RD7DOWNTO0_intermed_1 <= RIN.X.CTRL.RD ( 7 DOWNTO 0 );
		RIN_M_CTRL_RD7DOWNTO0_intermed_1 <= RIN.M.CTRL.RD ( 7 DOWNTO 0 );
		RIN_M_CTRL_RD7DOWNTO0_intermed_2 <= RIN_M_CTRL_RD7DOWNTO0_intermed_1;
		RIN_X_CTRL_TRAP_intermed_1 <= RIN.X.CTRL.TRAP;
		V_A_CTRL_TRAP_shadow_intermed_1 <= V_A_CTRL_TRAP_shadow;
		V_A_CTRL_TRAP_shadow_intermed_2 <= V_A_CTRL_TRAP_shadow_intermed_1;
		V_A_CTRL_TRAP_shadow_intermed_3 <= V_A_CTRL_TRAP_shadow_intermed_2;
		V_A_CTRL_TRAP_shadow_intermed_4 <= V_A_CTRL_TRAP_shadow_intermed_3;
		ICO_MEXC_intermed_1 <= ICO.MEXC;
		ICO_MEXC_intermed_2 <= ICO_MEXC_intermed_1;
		ICO_MEXC_intermed_3 <= ICO_MEXC_intermed_2;
		ICO_MEXC_intermed_4 <= ICO_MEXC_intermed_3;
		ICO_MEXC_intermed_5 <= ICO_MEXC_intermed_4;
		R_E_CTRL_TRAP_intermed_1 <= R.E.CTRL.TRAP;
		R_E_CTRL_TRAP_intermed_2 <= R_E_CTRL_TRAP_intermed_1;
		RIN_A_CTRL_TRAP_intermed_1 <= RIN.A.CTRL.TRAP;
		RIN_A_CTRL_TRAP_intermed_2 <= RIN_A_CTRL_TRAP_intermed_1;
		RIN_A_CTRL_TRAP_intermed_3 <= RIN_A_CTRL_TRAP_intermed_2;
		RIN_A_CTRL_TRAP_intermed_4 <= RIN_A_CTRL_TRAP_intermed_3;
		V_E_CTRL_TRAP_shadow_intermed_1 <= V_E_CTRL_TRAP_shadow;
		V_E_CTRL_TRAP_shadow_intermed_2 <= V_E_CTRL_TRAP_shadow_intermed_1;
		V_E_CTRL_TRAP_shadow_intermed_3 <= V_E_CTRL_TRAP_shadow_intermed_2;
		RIN_E_CTRL_TRAP_intermed_1 <= RIN.E.CTRL.TRAP;
		RIN_E_CTRL_TRAP_intermed_2 <= RIN_E_CTRL_TRAP_intermed_1;
		RIN_E_CTRL_TRAP_intermed_3 <= RIN_E_CTRL_TRAP_intermed_2;
		R_D_MEXC_intermed_1 <= R.D.MEXC;
		R_D_MEXC_intermed_2 <= R_D_MEXC_intermed_1;
		R_D_MEXC_intermed_3 <= R_D_MEXC_intermed_2;
		R_D_MEXC_intermed_4 <= R_D_MEXC_intermed_3;
		V_M_CTRL_TRAP_shadow_intermed_1 <= V_M_CTRL_TRAP_shadow;
		V_M_CTRL_TRAP_shadow_intermed_2 <= V_M_CTRL_TRAP_shadow_intermed_1;
		V_D_MEXC_shadow_intermed_1 <= V_D_MEXC_shadow;
		V_D_MEXC_shadow_intermed_2 <= V_D_MEXC_shadow_intermed_1;
		V_D_MEXC_shadow_intermed_3 <= V_D_MEXC_shadow_intermed_2;
		V_D_MEXC_shadow_intermed_4 <= V_D_MEXC_shadow_intermed_3;
		V_D_MEXC_shadow_intermed_5 <= V_D_MEXC_shadow_intermed_4;
		R_A_CTRL_TRAP_intermed_1 <= R.A.CTRL.TRAP;
		R_A_CTRL_TRAP_intermed_2 <= R_A_CTRL_TRAP_intermed_1;
		R_A_CTRL_TRAP_intermed_3 <= R_A_CTRL_TRAP_intermed_2;
		RIN_M_CTRL_TRAP_intermed_1 <= RIN.M.CTRL.TRAP;
		RIN_M_CTRL_TRAP_intermed_2 <= RIN_M_CTRL_TRAP_intermed_1;
		R_M_CTRL_TRAP_intermed_1 <= R.M.CTRL.TRAP;
		RIN_D_MEXC_intermed_1 <= RIN.D.MEXC;
		RIN_D_MEXC_intermed_2 <= RIN_D_MEXC_intermed_1;
		RIN_D_MEXC_intermed_3 <= RIN_D_MEXC_intermed_2;
		RIN_D_MEXC_intermed_4 <= RIN_D_MEXC_intermed_3;
		RIN_D_MEXC_intermed_5 <= RIN_D_MEXC_intermed_4;
		RIN_X_RESULT6DOWNTO0_intermed_1 <= RIN.X.RESULT ( 6 DOWNTO 0 );
		V_X_RESULT6DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO0_shadow;
		V_X_RESULT6DOWNTO0_shadow_intermed_2 <= V_X_RESULT6DOWNTO0_shadow_intermed_1;
		RIN_X_RESULT6DOWNTO0_intermed_1 <= RIN.X.RESULT( 6 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO0_intermed_2 <= RIN_X_RESULT6DOWNTO0_intermed_1;
		R_X_RESULT6DOWNTO0_intermed_1 <= R.X.RESULT( 6 DOWNTO 0 );
		RIN_D_PC_intermed_1 <= RIN.D.PC;
		RIN_D_PC_intermed_2 <= RIN_D_PC_intermed_1;
		RIN_D_PC_intermed_3 <= RIN_D_PC_intermed_2;
		RIN_D_PC_intermed_4 <= RIN_D_PC_intermed_3;
		RIN_D_PC_intermed_5 <= RIN_D_PC_intermed_4;
		RIN_A_CTRL_PC_intermed_1 <= RIN.A.CTRL.PC;
		RIN_A_CTRL_PC_intermed_2 <= RIN_A_CTRL_PC_intermed_1;
		RIN_A_CTRL_PC_intermed_3 <= RIN_A_CTRL_PC_intermed_2;
		RIN_A_CTRL_PC_intermed_4 <= RIN_A_CTRL_PC_intermed_3;
		R_A_CTRL_PC_intermed_1 <= R.A.CTRL.PC;
		R_A_CTRL_PC_intermed_2 <= R_A_CTRL_PC_intermed_1;
		R_A_CTRL_PC_intermed_3 <= R_A_CTRL_PC_intermed_2;
		V_E_CTRL_PC_shadow_intermed_1 <= V_E_CTRL_PC_shadow;
		V_E_CTRL_PC_shadow_intermed_2 <= V_E_CTRL_PC_shadow_intermed_1;
		V_E_CTRL_PC_shadow_intermed_3 <= V_E_CTRL_PC_shadow_intermed_2;
		R_M_CTRL_PC_intermed_1 <= R.M.CTRL.PC;
		R_E_CTRL_PC_intermed_1 <= R.E.CTRL.PC;
		R_E_CTRL_PC_intermed_2 <= R_E_CTRL_PC_intermed_1;
		RIN_M_CTRL_PC_intermed_1 <= RIN.M.CTRL.PC;
		RIN_M_CTRL_PC_intermed_2 <= RIN_M_CTRL_PC_intermed_1;
		V_M_CTRL_PC_shadow_intermed_1 <= V_M_CTRL_PC_shadow;
		V_M_CTRL_PC_shadow_intermed_2 <= V_M_CTRL_PC_shadow_intermed_1;
		V_A_CTRL_PC_shadow_intermed_1 <= V_A_CTRL_PC_shadow;
		V_A_CTRL_PC_shadow_intermed_2 <= V_A_CTRL_PC_shadow_intermed_1;
		V_A_CTRL_PC_shadow_intermed_3 <= V_A_CTRL_PC_shadow_intermed_2;
		V_A_CTRL_PC_shadow_intermed_4 <= V_A_CTRL_PC_shadow_intermed_3;
		R_D_PC_intermed_1 <= R.D.PC;
		R_D_PC_intermed_2 <= R_D_PC_intermed_1;
		R_D_PC_intermed_3 <= R_D_PC_intermed_2;
		R_D_PC_intermed_4 <= R_D_PC_intermed_3;
		RIN_E_CTRL_PC_intermed_1 <= RIN.E.CTRL.PC;
		RIN_E_CTRL_PC_intermed_2 <= RIN_E_CTRL_PC_intermed_1;
		RIN_E_CTRL_PC_intermed_3 <= RIN_E_CTRL_PC_intermed_2;
		RIN_X_CTRL_PC_intermed_1 <= RIN.X.CTRL.PC;
		V_D_PC_shadow_intermed_1 <= V_D_PC_shadow;
		V_D_PC_shadow_intermed_2 <= V_D_PC_shadow_intermed_1;
		V_D_PC_shadow_intermed_3 <= V_D_PC_shadow_intermed_2;
		V_D_PC_shadow_intermed_4 <= V_D_PC_shadow_intermed_3;
		V_D_PC_shadow_intermed_5 <= V_D_PC_shadow_intermed_4;
		RIN_A_CTRL_ANNUL_intermed_1 <= RIN.A.CTRL.ANNUL;
		RIN_A_CTRL_ANNUL_intermed_2 <= RIN_A_CTRL_ANNUL_intermed_1;
		RIN_A_CTRL_ANNUL_intermed_3 <= RIN_A_CTRL_ANNUL_intermed_2;
		RIN_A_CTRL_ANNUL_intermed_4 <= RIN_A_CTRL_ANNUL_intermed_3;
		RIN_A_CTRL_ANNUL_intermed_5 <= RIN_A_CTRL_ANNUL_intermed_4;
		R_A_CTRL_ANNUL_intermed_1 <= R.A.CTRL.ANNUL;
		R_A_CTRL_ANNUL_intermed_2 <= R_A_CTRL_ANNUL_intermed_1;
		R_A_CTRL_ANNUL_intermed_3 <= R_A_CTRL_ANNUL_intermed_2;
		R_A_CTRL_ANNUL_intermed_4 <= R_A_CTRL_ANNUL_intermed_3;
		R_X_ANNUL_ALL_intermed_1 <= R.X.ANNUL_ALL;
		R_X_ANNUL_ALL_intermed_2 <= R_X_ANNUL_ALL_intermed_1;
		R_X_ANNUL_ALL_intermed_3 <= R_X_ANNUL_ALL_intermed_2;
		R_X_ANNUL_ALL_intermed_4 <= R_X_ANNUL_ALL_intermed_3;
		RIN_X_CTRL_WREG_intermed_1 <= RIN.X.CTRL.WREG;
		RIN_M_CTRL_WREG_intermed_1 <= RIN.M.CTRL.WREG;
		RIN_M_CTRL_WREG_intermed_2 <= RIN_M_CTRL_WREG_intermed_1;
		RIN_A_CTRL_WREG_intermed_1 <= RIN.A.CTRL.WREG;
		RIN_A_CTRL_WREG_intermed_2 <= RIN_A_CTRL_WREG_intermed_1;
		RIN_A_CTRL_WREG_intermed_3 <= RIN_A_CTRL_WREG_intermed_2;
		RIN_A_CTRL_WREG_intermed_4 <= RIN_A_CTRL_WREG_intermed_3;
		V_A_CTRL_WREG_shadow_intermed_1 <= V_A_CTRL_WREG_shadow;
		V_A_CTRL_WREG_shadow_intermed_2 <= V_A_CTRL_WREG_shadow_intermed_1;
		V_A_CTRL_WREG_shadow_intermed_3 <= V_A_CTRL_WREG_shadow_intermed_2;
		V_A_CTRL_WREG_shadow_intermed_4 <= V_A_CTRL_WREG_shadow_intermed_3;
		R_A_CTRL_WREG_intermed_1 <= R.A.CTRL.WREG;
		R_A_CTRL_WREG_intermed_2 <= R_A_CTRL_WREG_intermed_1;
		R_A_CTRL_WREG_intermed_3 <= R_A_CTRL_WREG_intermed_2;
		V_X_ANNUL_ALL_shadow_intermed_1 <= V_X_ANNUL_ALL_shadow;
		V_X_ANNUL_ALL_shadow_intermed_2 <= V_X_ANNUL_ALL_shadow_intermed_1;
		V_X_ANNUL_ALL_shadow_intermed_3 <= V_X_ANNUL_ALL_shadow_intermed_2;
		V_X_ANNUL_ALL_shadow_intermed_4 <= V_X_ANNUL_ALL_shadow_intermed_3;
		R_M_CTRL_WREG_intermed_1 <= R.M.CTRL.WREG;
		RIN_X_ANNUL_ALL_intermed_1 <= RIN.X.ANNUL_ALL;
		RIN_X_ANNUL_ALL_intermed_2 <= RIN_X_ANNUL_ALL_intermed_1;
		RIN_X_ANNUL_ALL_intermed_3 <= RIN_X_ANNUL_ALL_intermed_2;
		RIN_X_ANNUL_ALL_intermed_4 <= RIN_X_ANNUL_ALL_intermed_3;
		RIN_X_ANNUL_ALL_intermed_5 <= RIN_X_ANNUL_ALL_intermed_4;
		V_M_CTRL_WREG_shadow_intermed_1 <= V_M_CTRL_WREG_shadow;
		V_M_CTRL_WREG_shadow_intermed_2 <= V_M_CTRL_WREG_shadow_intermed_1;
		R_E_CTRL_WREG_intermed_1 <= R.E.CTRL.WREG;
		R_E_CTRL_WREG_intermed_2 <= R_E_CTRL_WREG_intermed_1;
		V_A_CTRL_ANNUL_shadow_intermed_1 <= V_A_CTRL_ANNUL_shadow;
		V_A_CTRL_ANNUL_shadow_intermed_2 <= V_A_CTRL_ANNUL_shadow_intermed_1;
		V_A_CTRL_ANNUL_shadow_intermed_3 <= V_A_CTRL_ANNUL_shadow_intermed_2;
		V_A_CTRL_ANNUL_shadow_intermed_4 <= V_A_CTRL_ANNUL_shadow_intermed_3;
		RIN_E_CTRL_WREG_intermed_1 <= RIN.E.CTRL.WREG;
		RIN_E_CTRL_WREG_intermed_2 <= RIN_E_CTRL_WREG_intermed_1;
		RIN_E_CTRL_WREG_intermed_3 <= RIN_E_CTRL_WREG_intermed_2;
		V_E_CTRL_WREG_shadow_intermed_1 <= V_E_CTRL_WREG_shadow;
		V_E_CTRL_WREG_shadow_intermed_2 <= V_E_CTRL_WREG_shadow_intermed_1;
		V_E_CTRL_WREG_shadow_intermed_3 <= V_E_CTRL_WREG_shadow_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_3 <= RIN_M_CTRL_PC31DOWNTO2_intermed_2;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC ( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_5 <= V_D_PC31DOWNTO2_shadow_intermed_4;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_5 <= RIN_D_PC31DOWNTO2_intermed_4;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC ( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC ( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC ( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_2 <= RIN_X_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC ( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		R_D_PC31DOWNTO2_intermed_4 <= R_D_PC31DOWNTO2_intermed_3;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC ( 31 DOWNTO 2 );
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 2 );
		R_M_CTRL_PC31DOWNTO2_intermed_2 <= R_M_CTRL_PC31DOWNTO2_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		RIN_A_CTRL_PC31DOWNTO2_intermed_5 <= RIN_A_CTRL_PC31DOWNTO2_intermed_4;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_4 <= R_A_CTRL_PC31DOWNTO2_intermed_3;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC ( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		R_X_CTRL_PC31DOWNTO2_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 2 );
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_3 <= R_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_4 <= RIN_E_CTRL_PC31DOWNTO2_intermed_3;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO2_shadow;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_5 <= V_D_PC31DOWNTO2_shadow_intermed_4;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_5 <= RIN_D_PC31DOWNTO2_intermed_4;
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 2 );
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		R_D_PC31DOWNTO2_intermed_4 <= R_D_PC31DOWNTO2_intermed_3;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 2 );
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		V_X_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_X_CTRL_TT3DOWNTO0_shadow;
		V_X_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_X_CTRL_TT3DOWNTO0_shadow_intermed_1;
		R_M_CTRL_TT3DOWNTO0_intermed_1 <= R.M.CTRL.TT( 3 DOWNTO 0 );
		R_M_CTRL_TT3DOWNTO0_intermed_2 <= R_M_CTRL_TT3DOWNTO0_intermed_1;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_3 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2;
		R_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= R.X.RESULT( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		R_X_RESULT6DOWNTO03DOWNTO0_intermed_2 <= R_X_RESULT6DOWNTO03DOWNTO0_intermed_1;
		R_A_CTRL_TT3DOWNTO0_intermed_1 <= R.A.CTRL.TT( 3 DOWNTO 0 );
		R_A_CTRL_TT3DOWNTO0_intermed_2 <= R_A_CTRL_TT3DOWNTO0_intermed_1;
		R_A_CTRL_TT3DOWNTO0_intermed_3 <= R_A_CTRL_TT3DOWNTO0_intermed_2;
		R_A_CTRL_TT3DOWNTO0_intermed_4 <= R_A_CTRL_TT3DOWNTO0_intermed_3;
		RIN_A_CTRL_TT3DOWNTO0_intermed_1 <= RIN.A.CTRL.TT( 3 DOWNTO 0 );
		RIN_A_CTRL_TT3DOWNTO0_intermed_2 <= RIN_A_CTRL_TT3DOWNTO0_intermed_1;
		RIN_A_CTRL_TT3DOWNTO0_intermed_3 <= RIN_A_CTRL_TT3DOWNTO0_intermed_2;
		RIN_A_CTRL_TT3DOWNTO0_intermed_4 <= RIN_A_CTRL_TT3DOWNTO0_intermed_3;
		RIN_A_CTRL_TT3DOWNTO0_intermed_5 <= RIN_A_CTRL_TT3DOWNTO0_intermed_4;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_A_CTRL_TT3DOWNTO0_shadow;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_1;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_3 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_2;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_4 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_3;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_5 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_4;
		RIN_W_S_TT3DOWNTO0_intermed_1 <= RIN.W.S.TT( 3 DOWNTO 0 );
		RIN_W_S_TT3DOWNTO0_intermed_2 <= RIN_W_S_TT3DOWNTO0_intermed_1;
		R_E_CTRL_TT3DOWNTO0_intermed_1 <= R.E.CTRL.TT( 3 DOWNTO 0 );
		R_E_CTRL_TT3DOWNTO0_intermed_2 <= R_E_CTRL_TT3DOWNTO0_intermed_1;
		R_E_CTRL_TT3DOWNTO0_intermed_3 <= R_E_CTRL_TT3DOWNTO0_intermed_2;
		RIN_W_S_TT3DOWNTO0_intermed_1 <= RIN.W.S.TT ( 3 DOWNTO 0 );
		RIN_M_CTRL_TT3DOWNTO0_intermed_1 <= RIN.M.CTRL.TT( 3 DOWNTO 0 );
		RIN_M_CTRL_TT3DOWNTO0_intermed_2 <= RIN_M_CTRL_TT3DOWNTO0_intermed_1;
		RIN_M_CTRL_TT3DOWNTO0_intermed_3 <= RIN_M_CTRL_TT3DOWNTO0_intermed_2;
		V_M_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_M_CTRL_TT3DOWNTO0_shadow;
		V_M_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_M_CTRL_TT3DOWNTO0_shadow_intermed_1;
		V_M_CTRL_TT3DOWNTO0_shadow_intermed_3 <= V_M_CTRL_TT3DOWNTO0_shadow_intermed_2;
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= RIN.X.RESULT( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2 <= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1;
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_3 <= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2;
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= RIN.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2 <= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1;
		R_W_S_TT3DOWNTO0_intermed_1 <= R.W.S.TT( 3 DOWNTO 0 );
		R_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= R.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_E_CTRL_TT3DOWNTO0_shadow;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_E_CTRL_TT3DOWNTO0_shadow_intermed_1;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_3 <= V_E_CTRL_TT3DOWNTO0_shadow_intermed_2;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_4 <= V_E_CTRL_TT3DOWNTO0_shadow_intermed_3;
		RIN_X_CTRL_TT3DOWNTO0_intermed_1 <= RIN.X.CTRL.TT( 3 DOWNTO 0 );
		RIN_X_CTRL_TT3DOWNTO0_intermed_2 <= RIN_X_CTRL_TT3DOWNTO0_intermed_1;
		V_W_S_TT3DOWNTO0_shadow_intermed_1 <= V_W_S_TT3DOWNTO0_shadow;
		V_W_S_TT3DOWNTO0_shadow_intermed_2 <= V_W_S_TT3DOWNTO0_shadow_intermed_1;
		R_X_CTRL_TT3DOWNTO0_intermed_1 <= R.X.CTRL.TT( 3 DOWNTO 0 );
		RIN_E_CTRL_TT3DOWNTO0_intermed_1 <= RIN.E.CTRL.TT( 3 DOWNTO 0 );
		RIN_E_CTRL_TT3DOWNTO0_intermed_2 <= RIN_E_CTRL_TT3DOWNTO0_intermed_1;
		RIN_E_CTRL_TT3DOWNTO0_intermed_3 <= RIN_E_CTRL_TT3DOWNTO0_intermed_2;
		RIN_E_CTRL_TT3DOWNTO0_intermed_4 <= RIN_E_CTRL_TT3DOWNTO0_intermed_3;
		XC_VECTT3DOWNTO0_shadow_intermed_1 <= XC_VECTT3DOWNTO0_shadow;
		V_M_RESULT1DOWNTO0_shadow_intermed_1 <= V_M_RESULT1DOWNTO0_shadow;
		V_M_RESULT1DOWNTO0_shadow_intermed_2 <= V_M_RESULT1DOWNTO0_shadow_intermed_1;
		RIN_M_RESULT1DOWNTO0_intermed_1 <= RIN.M.RESULT( 1 DOWNTO 0 );
		RIN_M_RESULT1DOWNTO0_intermed_2 <= RIN_M_RESULT1DOWNTO0_intermed_1;
		R_M_RESULT1DOWNTO0_intermed_1 <= R.M.RESULT( 1 DOWNTO 0 );
		RIN_M_RESULT1DOWNTO0_intermed_1 <= RIN.M.RESULT ( 1 DOWNTO 0 );
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA ( 0 )( 31 );
		RIN_X_DATA031_intermed_2 <= RIN_X_DATA031_intermed_1;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_2 <= V_X_DATA031_shadow_intermed_1;
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_2 <= V_X_DATA031_shadow_intermed_1;
		V_X_DATA031_shadow_intermed_3 <= V_X_DATA031_shadow_intermed_2;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA( 0 )( 31 );
		RIN_X_DATA031_intermed_2 <= RIN_X_DATA031_intermed_1;
		RIN_X_DATA031_intermed_3 <= RIN_X_DATA031_intermed_2;
		DCO_DATA031_intermed_1 <= DCO.DATA ( 0 )( 31 );
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA ( 0 ) ( 31 );
		R_X_DATA031_intermed_1 <= R.X.DATA( 0 )( 31 );
		R_X_DATA031_intermed_2 <= R_X_DATA031_intermed_1;
		R_X_DATA031_intermed_1 <= R.X.DATA ( 0 )( 31 );
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA ( 0 )( 31 );
		V_X_DATA031_shadow_intermed_1 <= V_X_DATA031_shadow;
		V_X_DATA031_shadow_intermed_2 <= V_X_DATA031_shadow_intermed_1;
		RIN_X_DATA031_intermed_1 <= RIN.X.DATA( 0 )( 31 );
		RIN_X_DATA031_intermed_2 <= RIN_X_DATA031_intermed_1;
		DCO_DATA031_intermed_1 <= DCO.DATA ( 0 )( 31 );
		R_X_DATA031_intermed_1 <= R.X.DATA( 0 )( 31 );
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		V_A_CTRL_INST19_shadow_intermed_3 <= V_A_CTRL_INST19_shadow_intermed_2;
		V_E_CTRL_INST19_shadow_intermed_1 <= V_E_CTRL_INST19_shadow;
		V_E_CTRL_INST19_shadow_intermed_2 <= V_E_CTRL_INST19_shadow_intermed_1;
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST ( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		RIN_A_CTRL_INST19_intermed_3 <= RIN_A_CTRL_INST19_intermed_2;
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST ( 19 );
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST( 19 );
		RIN_E_CTRL_INST19_intermed_2 <= RIN_E_CTRL_INST19_intermed_1;
		DE_INST19_shadow_intermed_1 <= DE_INST19_shadow;
		DE_INST19_shadow_intermed_2 <= DE_INST19_shadow_intermed_1;
		R_E_CTRL_INST19_intermed_1 <= R.E.CTRL.INST( 19 );
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST( 19 );
		R_A_CTRL_INST19_intermed_2 <= R_A_CTRL_INST19_intermed_1;
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST ( 19 );
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		RIN_A_CTRL_INST20_intermed_1 <= RIN.A.CTRL.INST ( 20 );
		RIN_A_CTRL_INST20_intermed_2 <= RIN_A_CTRL_INST20_intermed_1;
		R_A_CTRL_INST20_intermed_1 <= R.A.CTRL.INST ( 20 );
		RIN_A_CTRL_INST20_intermed_1 <= RIN.A.CTRL.INST( 20 );
		RIN_A_CTRL_INST20_intermed_2 <= RIN_A_CTRL_INST20_intermed_1;
		RIN_A_CTRL_INST20_intermed_3 <= RIN_A_CTRL_INST20_intermed_2;
		V_E_CTRL_INST20_shadow_intermed_1 <= V_E_CTRL_INST20_shadow;
		V_E_CTRL_INST20_shadow_intermed_2 <= V_E_CTRL_INST20_shadow_intermed_1;
		V_A_CTRL_INST20_shadow_intermed_1 <= V_A_CTRL_INST20_shadow;
		V_A_CTRL_INST20_shadow_intermed_2 <= V_A_CTRL_INST20_shadow_intermed_1;
		V_A_CTRL_INST20_shadow_intermed_3 <= V_A_CTRL_INST20_shadow_intermed_2;
		RIN_E_CTRL_INST20_intermed_1 <= RIN.E.CTRL.INST( 20 );
		RIN_E_CTRL_INST20_intermed_2 <= RIN_E_CTRL_INST20_intermed_1;
		V_A_CTRL_INST20_shadow_intermed_1 <= V_A_CTRL_INST20_shadow;
		V_A_CTRL_INST20_shadow_intermed_2 <= V_A_CTRL_INST20_shadow_intermed_1;
		RIN_E_CTRL_INST20_intermed_1 <= RIN.E.CTRL.INST ( 20 );
		R_E_CTRL_INST20_intermed_1 <= R.E.CTRL.INST( 20 );
		DE_INST20_shadow_intermed_1 <= DE_INST20_shadow;
		DE_INST20_shadow_intermed_2 <= DE_INST20_shadow_intermed_1;
		R_A_CTRL_INST20_intermed_1 <= R.A.CTRL.INST( 20 );
		R_A_CTRL_INST20_intermed_2 <= R_A_CTRL_INST20_intermed_1;
		V_X_DATA00_shadow_intermed_1 <= V_X_DATA00_shadow;
		V_X_DATA00_shadow_intermed_2 <= V_X_DATA00_shadow_intermed_1;
		RIN_X_DATA00_intermed_1 <= RIN.X.DATA ( 0 ) ( 0 );
		R_X_DATA00_intermed_1 <= R.X.DATA( 0 )( 0 );
		R_X_DATA00_intermed_2 <= R_X_DATA00_intermed_1;
		RIN_X_DATA00_intermed_1 <= RIN.X.DATA ( 0 )( 0 );
		RIN_X_DATA00_intermed_2 <= RIN_X_DATA00_intermed_1;
		DCO_DATA00_intermed_1 <= DCO.DATA ( 0 )( 0 );
		V_X_DATA00_shadow_intermed_1 <= V_X_DATA00_shadow;
		V_X_DATA00_shadow_intermed_2 <= V_X_DATA00_shadow_intermed_1;
		V_X_DATA00_shadow_intermed_3 <= V_X_DATA00_shadow_intermed_2;
		R_X_DATA00_intermed_1 <= R.X.DATA ( 0 )( 0 );
		RIN_X_DATA00_intermed_1 <= RIN.X.DATA( 0 )( 0 );
		RIN_X_DATA00_intermed_2 <= RIN_X_DATA00_intermed_1;
		RIN_X_DATA00_intermed_3 <= RIN_X_DATA00_intermed_2;
		R_X_DATA00_intermed_1 <= R.X.DATA( 0 )( 0 );
		RIN_X_DATA00_intermed_1 <= RIN.X.DATA ( 0 )( 0 );
		DCO_DATA00_intermed_1 <= DCO.DATA ( 0 )( 0 );
		V_X_DATA00_shadow_intermed_1 <= V_X_DATA00_shadow;
		V_X_DATA00_shadow_intermed_2 <= V_X_DATA00_shadow_intermed_1;
		RIN_X_DATA00_intermed_1 <= RIN.X.DATA( 0 )( 0 );
		RIN_X_DATA00_intermed_2 <= RIN_X_DATA00_intermed_1;
		RIN_X_DATA04DOWNTO0_intermed_1 <= RIN.X.DATA ( 0 ) ( 4 DOWNTO 0 );
		R_X_DATA04DOWNTO0_intermed_1 <= R.X.DATA( 0 )( 4 DOWNTO 0 );
		R_X_DATA04DOWNTO0_intermed_2 <= R_X_DATA04DOWNTO0_intermed_1;
		R_X_DATA04DOWNTO0_intermed_1 <= R.X.DATA ( 0 )( 4 DOWNTO 0 );
		RIN_X_DATA04DOWNTO0_intermed_1 <= RIN.X.DATA( 0 )( 4 DOWNTO 0 );
		RIN_X_DATA04DOWNTO0_intermed_2 <= RIN_X_DATA04DOWNTO0_intermed_1;
		RIN_X_DATA04DOWNTO0_intermed_3 <= RIN_X_DATA04DOWNTO0_intermed_2;
		V_X_DATA04DOWNTO0_shadow_intermed_1 <= V_X_DATA04DOWNTO0_shadow;
		V_X_DATA04DOWNTO0_shadow_intermed_2 <= V_X_DATA04DOWNTO0_shadow_intermed_1;
		V_X_DATA04DOWNTO0_shadow_intermed_1 <= V_X_DATA04DOWNTO0_shadow;
		V_X_DATA04DOWNTO0_shadow_intermed_2 <= V_X_DATA04DOWNTO0_shadow_intermed_1;
		V_X_DATA04DOWNTO0_shadow_intermed_3 <= V_X_DATA04DOWNTO0_shadow_intermed_2;
		RIN_X_DATA04DOWNTO0_intermed_1 <= RIN.X.DATA ( 0 )( 4 DOWNTO 0 );
		RIN_X_DATA04DOWNTO0_intermed_2 <= RIN_X_DATA04DOWNTO0_intermed_1;
		DCO_DATA04DOWNTO0_intermed_1 <= DCO.DATA ( 0 )( 4 DOWNTO 0 );
		R_X_DATA04DOWNTO0_intermed_1 <= R.X.DATA( 0 )( 4 DOWNTO 0 );
		RIN_X_DATA04DOWNTO0_intermed_1 <= RIN.X.DATA( 0 )( 4 DOWNTO 0 );
		RIN_X_DATA04DOWNTO0_intermed_2 <= RIN_X_DATA04DOWNTO0_intermed_1;
		V_X_DATA04DOWNTO0_shadow_intermed_1 <= V_X_DATA04DOWNTO0_shadow;
		V_X_DATA04DOWNTO0_shadow_intermed_2 <= V_X_DATA04DOWNTO0_shadow_intermed_1;
		DCO_DATA04DOWNTO0_intermed_1 <= DCO.DATA ( 0 )( 4 DOWNTO 0 );
		RIN_X_DATA04DOWNTO0_intermed_1 <= RIN.X.DATA ( 0 )( 4 DOWNTO 0 );
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC ( 31 DOWNTO 2 );
		R_A_CTRL_INST24_intermed_1 <= R.A.CTRL.INST( 24 );
		R_A_CTRL_INST24_intermed_2 <= R_A_CTRL_INST24_intermed_1;
		RIN_E_CTRL_INST24_intermed_1 <= RIN.E.CTRL.INST( 24 );
		RIN_E_CTRL_INST24_intermed_2 <= RIN_E_CTRL_INST24_intermed_1;
		RIN_A_CTRL_INST24_intermed_1 <= RIN.A.CTRL.INST( 24 );
		RIN_A_CTRL_INST24_intermed_2 <= RIN_A_CTRL_INST24_intermed_1;
		RIN_A_CTRL_INST24_intermed_3 <= RIN_A_CTRL_INST24_intermed_2;
		R_E_CTRL_INST24_intermed_1 <= R.E.CTRL.INST( 24 );
		R_A_CTRL_INST24_intermed_1 <= R.A.CTRL.INST ( 24 );
		V_A_CTRL_INST24_shadow_intermed_1 <= V_A_CTRL_INST24_shadow;
		V_A_CTRL_INST24_shadow_intermed_2 <= V_A_CTRL_INST24_shadow_intermed_1;
		V_A_CTRL_INST24_shadow_intermed_3 <= V_A_CTRL_INST24_shadow_intermed_2;
		V_E_CTRL_INST24_shadow_intermed_1 <= V_E_CTRL_INST24_shadow;
		V_E_CTRL_INST24_shadow_intermed_2 <= V_E_CTRL_INST24_shadow_intermed_1;
		DE_INST24_shadow_intermed_1 <= DE_INST24_shadow;
		DE_INST24_shadow_intermed_2 <= DE_INST24_shadow_intermed_1;
		RIN_A_CTRL_INST24_intermed_1 <= RIN.A.CTRL.INST ( 24 );
		RIN_A_CTRL_INST24_intermed_2 <= RIN_A_CTRL_INST24_intermed_1;
		V_A_CTRL_INST24_shadow_intermed_1 <= V_A_CTRL_INST24_shadow;
		V_A_CTRL_INST24_shadow_intermed_2 <= V_A_CTRL_INST24_shadow_intermed_1;
		RIN_E_CTRL_INST24_intermed_1 <= RIN.E.CTRL.INST ( 24 );
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST ( 19 );
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		DE_INST19_shadow_intermed_1 <= DE_INST19_shadow;
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST( 19 );
		RIN_M_Y31_intermed_1 <= RIN.M.Y ( 31 );
		V_M_Y31_shadow_intermed_1 <= V_M_Y31_shadow;
		V_M_Y31_shadow_intermed_2 <= V_M_Y31_shadow_intermed_1;
		RIN_M_Y31_intermed_1 <= RIN.M.Y( 31 );
		RIN_M_Y31_intermed_2 <= RIN_M_Y31_intermed_1;
		R_M_Y31_intermed_1 <= R.M.Y( 31 );
		DSUIN_CRDY2_intermed_1 <= DSUIN.CRDY ( 2 );
		VDSU_CRDY2_shadow_intermed_1 <= VDSU_CRDY2_shadow;
		VDSU_CRDY2_shadow_intermed_2 <= VDSU_CRDY2_shadow_intermed_1;
		DSUIN_CRDY2_intermed_1 <= DSUIN.CRDY( 2 );
		DSUIN_CRDY2_intermed_2 <= DSUIN_CRDY2_intermed_1;
		DSUR_CRDY2_intermed_1 <= DSUR.CRDY( 2 );
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC ( 31 DOWNTO 2 );
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC ( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC ( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC ( 31 DOWNTO 2 );
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		DE_INST_shadow_intermed_1 <= DE_INST_shadow;
		DE_INST_shadow_intermed_2 <= DE_INST_shadow_intermed_1;
		V_A_CTRL_INST_shadow_intermed_1 <= V_A_CTRL_INST_shadow;
		V_A_CTRL_INST_shadow_intermed_2 <= V_A_CTRL_INST_shadow_intermed_1;
		RIN_A_CTRL_INST_intermed_1 <= RIN.A.CTRL.INST;
		RIN_A_CTRL_INST_intermed_2 <= RIN_A_CTRL_INST_intermed_1;
		RIN_E_CTRL_INST_intermed_1 <= RIN.E.CTRL.INST;
		R_A_CTRL_INST_intermed_1 <= R.A.CTRL.INST;
		RIN_D_CNT_intermed_1 <= RIN.D.CNT;
		RIN_D_CNT_intermed_2 <= RIN_D_CNT_intermed_1;
		RIN_D_CNT_intermed_3 <= RIN_D_CNT_intermed_2;
		V_A_CTRL_CNT_shadow_intermed_1 <= V_A_CTRL_CNT_shadow;
		V_A_CTRL_CNT_shadow_intermed_2 <= V_A_CTRL_CNT_shadow_intermed_1;
		R_A_CTRL_CNT_intermed_1 <= R.A.CTRL.CNT;
		V_D_CNT_shadow_intermed_1 <= V_D_CNT_shadow;
		V_D_CNT_shadow_intermed_2 <= V_D_CNT_shadow_intermed_1;
		V_D_CNT_shadow_intermed_3 <= V_D_CNT_shadow_intermed_2;
		R_D_CNT_intermed_1 <= R.D.CNT;
		R_D_CNT_intermed_2 <= R_D_CNT_intermed_1;
		RIN_A_CTRL_CNT_intermed_1 <= RIN.A.CTRL.CNT;
		RIN_A_CTRL_CNT_intermed_2 <= RIN_A_CTRL_CNT_intermed_1;
		RIN_E_CTRL_CNT_intermed_1 <= RIN.E.CTRL.CNT;
		V_A_CTRL_TRAP_shadow_intermed_1 <= V_A_CTRL_TRAP_shadow;
		V_A_CTRL_TRAP_shadow_intermed_2 <= V_A_CTRL_TRAP_shadow_intermed_1;
		ICO_MEXC_intermed_1 <= ICO.MEXC;
		ICO_MEXC_intermed_2 <= ICO_MEXC_intermed_1;
		ICO_MEXC_intermed_3 <= ICO_MEXC_intermed_2;
		RIN_A_CTRL_TRAP_intermed_1 <= RIN.A.CTRL.TRAP;
		RIN_A_CTRL_TRAP_intermed_2 <= RIN_A_CTRL_TRAP_intermed_1;
		RIN_E_CTRL_TRAP_intermed_1 <= RIN.E.CTRL.TRAP;
		R_D_MEXC_intermed_1 <= R.D.MEXC;
		R_D_MEXC_intermed_2 <= R_D_MEXC_intermed_1;
		V_D_MEXC_shadow_intermed_1 <= V_D_MEXC_shadow;
		V_D_MEXC_shadow_intermed_2 <= V_D_MEXC_shadow_intermed_1;
		V_D_MEXC_shadow_intermed_3 <= V_D_MEXC_shadow_intermed_2;
		R_A_CTRL_TRAP_intermed_1 <= R.A.CTRL.TRAP;
		RIN_D_MEXC_intermed_1 <= RIN.D.MEXC;
		RIN_D_MEXC_intermed_2 <= RIN_D_MEXC_intermed_1;
		RIN_D_MEXC_intermed_3 <= RIN_D_MEXC_intermed_2;
		R_A_CTRL_PV_intermed_1 <= R.A.CTRL.PV;
		RIN_E_CTRL_PV_intermed_1 <= RIN.E.CTRL.PV;
		V_A_CTRL_PV_shadow_intermed_1 <= V_A_CTRL_PV_shadow;
		V_A_CTRL_PV_shadow_intermed_2 <= V_A_CTRL_PV_shadow_intermed_1;
		RIN_A_CTRL_PV_intermed_1 <= RIN.A.CTRL.PV;
		RIN_A_CTRL_PV_intermed_2 <= RIN_A_CTRL_PV_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC ( 31 DOWNTO 2 );
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC ( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC ( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC ( 31 DOWNTO 2 );
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 2 );
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC ( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		R_E_CTRL_INST_intermed_1 <= R.E.CTRL.INST;
		DE_INST_shadow_intermed_1 <= DE_INST_shadow;
		DE_INST_shadow_intermed_2 <= DE_INST_shadow_intermed_1;
		DE_INST_shadow_intermed_3 <= DE_INST_shadow_intermed_2;
		V_A_CTRL_INST_shadow_intermed_1 <= V_A_CTRL_INST_shadow;
		V_A_CTRL_INST_shadow_intermed_2 <= V_A_CTRL_INST_shadow_intermed_1;
		V_A_CTRL_INST_shadow_intermed_3 <= V_A_CTRL_INST_shadow_intermed_2;
		V_E_CTRL_INST_shadow_intermed_1 <= V_E_CTRL_INST_shadow;
		V_E_CTRL_INST_shadow_intermed_2 <= V_E_CTRL_INST_shadow_intermed_1;
		RIN_A_CTRL_INST_intermed_1 <= RIN.A.CTRL.INST;
		RIN_A_CTRL_INST_intermed_2 <= RIN_A_CTRL_INST_intermed_1;
		RIN_A_CTRL_INST_intermed_3 <= RIN_A_CTRL_INST_intermed_2;
		RIN_M_CTRL_INST_intermed_1 <= RIN.M.CTRL.INST;
		RIN_E_CTRL_INST_intermed_1 <= RIN.E.CTRL.INST;
		RIN_E_CTRL_INST_intermed_2 <= RIN_E_CTRL_INST_intermed_1;
		R_A_CTRL_INST_intermed_1 <= R.A.CTRL.INST;
		R_A_CTRL_INST_intermed_2 <= R_A_CTRL_INST_intermed_1;
		V_E_CTRL_CNT_shadow_intermed_1 <= V_E_CTRL_CNT_shadow;
		V_E_CTRL_CNT_shadow_intermed_2 <= V_E_CTRL_CNT_shadow_intermed_1;
		RIN_D_CNT_intermed_1 <= RIN.D.CNT;
		RIN_D_CNT_intermed_2 <= RIN_D_CNT_intermed_1;
		RIN_D_CNT_intermed_3 <= RIN_D_CNT_intermed_2;
		RIN_D_CNT_intermed_4 <= RIN_D_CNT_intermed_3;
		V_A_CTRL_CNT_shadow_intermed_1 <= V_A_CTRL_CNT_shadow;
		V_A_CTRL_CNT_shadow_intermed_2 <= V_A_CTRL_CNT_shadow_intermed_1;
		V_A_CTRL_CNT_shadow_intermed_3 <= V_A_CTRL_CNT_shadow_intermed_2;
		R_A_CTRL_CNT_intermed_1 <= R.A.CTRL.CNT;
		R_A_CTRL_CNT_intermed_2 <= R_A_CTRL_CNT_intermed_1;
		V_D_CNT_shadow_intermed_1 <= V_D_CNT_shadow;
		V_D_CNT_shadow_intermed_2 <= V_D_CNT_shadow_intermed_1;
		V_D_CNT_shadow_intermed_3 <= V_D_CNT_shadow_intermed_2;
		V_D_CNT_shadow_intermed_4 <= V_D_CNT_shadow_intermed_3;
		R_D_CNT_intermed_1 <= R.D.CNT;
		R_D_CNT_intermed_2 <= R_D_CNT_intermed_1;
		R_D_CNT_intermed_3 <= R_D_CNT_intermed_2;
		R_E_CTRL_CNT_intermed_1 <= R.E.CTRL.CNT;
		RIN_A_CTRL_CNT_intermed_1 <= RIN.A.CTRL.CNT;
		RIN_A_CTRL_CNT_intermed_2 <= RIN_A_CTRL_CNT_intermed_1;
		RIN_A_CTRL_CNT_intermed_3 <= RIN_A_CTRL_CNT_intermed_2;
		RIN_M_CTRL_CNT_intermed_1 <= RIN.M.CTRL.CNT;
		RIN_E_CTRL_CNT_intermed_1 <= RIN.E.CTRL.CNT;
		RIN_E_CTRL_CNT_intermed_2 <= RIN_E_CTRL_CNT_intermed_1;
		V_A_CTRL_TRAP_shadow_intermed_1 <= V_A_CTRL_TRAP_shadow;
		V_A_CTRL_TRAP_shadow_intermed_2 <= V_A_CTRL_TRAP_shadow_intermed_1;
		V_A_CTRL_TRAP_shadow_intermed_3 <= V_A_CTRL_TRAP_shadow_intermed_2;
		ICO_MEXC_intermed_1 <= ICO.MEXC;
		ICO_MEXC_intermed_2 <= ICO_MEXC_intermed_1;
		ICO_MEXC_intermed_3 <= ICO_MEXC_intermed_2;
		ICO_MEXC_intermed_4 <= ICO_MEXC_intermed_3;
		R_E_CTRL_TRAP_intermed_1 <= R.E.CTRL.TRAP;
		RIN_A_CTRL_TRAP_intermed_1 <= RIN.A.CTRL.TRAP;
		RIN_A_CTRL_TRAP_intermed_2 <= RIN_A_CTRL_TRAP_intermed_1;
		RIN_A_CTRL_TRAP_intermed_3 <= RIN_A_CTRL_TRAP_intermed_2;
		V_E_CTRL_TRAP_shadow_intermed_1 <= V_E_CTRL_TRAP_shadow;
		V_E_CTRL_TRAP_shadow_intermed_2 <= V_E_CTRL_TRAP_shadow_intermed_1;
		RIN_E_CTRL_TRAP_intermed_1 <= RIN.E.CTRL.TRAP;
		RIN_E_CTRL_TRAP_intermed_2 <= RIN_E_CTRL_TRAP_intermed_1;
		R_D_MEXC_intermed_1 <= R.D.MEXC;
		R_D_MEXC_intermed_2 <= R_D_MEXC_intermed_1;
		R_D_MEXC_intermed_3 <= R_D_MEXC_intermed_2;
		V_D_MEXC_shadow_intermed_1 <= V_D_MEXC_shadow;
		V_D_MEXC_shadow_intermed_2 <= V_D_MEXC_shadow_intermed_1;
		V_D_MEXC_shadow_intermed_3 <= V_D_MEXC_shadow_intermed_2;
		V_D_MEXC_shadow_intermed_4 <= V_D_MEXC_shadow_intermed_3;
		R_A_CTRL_TRAP_intermed_1 <= R.A.CTRL.TRAP;
		R_A_CTRL_TRAP_intermed_2 <= R_A_CTRL_TRAP_intermed_1;
		RIN_M_CTRL_TRAP_intermed_1 <= RIN.M.CTRL.TRAP;
		RIN_D_MEXC_intermed_1 <= RIN.D.MEXC;
		RIN_D_MEXC_intermed_2 <= RIN_D_MEXC_intermed_1;
		RIN_D_MEXC_intermed_3 <= RIN_D_MEXC_intermed_2;
		RIN_D_MEXC_intermed_4 <= RIN_D_MEXC_intermed_3;
		V_E_CTRL_PV_shadow_intermed_1 <= V_E_CTRL_PV_shadow;
		V_E_CTRL_PV_shadow_intermed_2 <= V_E_CTRL_PV_shadow_intermed_1;
		R_E_CTRL_PV_intermed_1 <= R.E.CTRL.PV;
		R_A_CTRL_PV_intermed_1 <= R.A.CTRL.PV;
		R_A_CTRL_PV_intermed_2 <= R_A_CTRL_PV_intermed_1;
		RIN_E_CTRL_PV_intermed_1 <= RIN.E.CTRL.PV;
		RIN_E_CTRL_PV_intermed_2 <= RIN_E_CTRL_PV_intermed_1;
		RIN_M_CTRL_PV_intermed_1 <= RIN.M.CTRL.PV;
		V_A_CTRL_PV_shadow_intermed_1 <= V_A_CTRL_PV_shadow;
		V_A_CTRL_PV_shadow_intermed_2 <= V_A_CTRL_PV_shadow_intermed_1;
		V_A_CTRL_PV_shadow_intermed_3 <= V_A_CTRL_PV_shadow_intermed_2;
		RIN_A_CTRL_PV_intermed_1 <= RIN.A.CTRL.PV;
		RIN_A_CTRL_PV_intermed_2 <= RIN_A_CTRL_PV_intermed_1;
		RIN_A_CTRL_PV_intermed_3 <= RIN_A_CTRL_PV_intermed_2;
		R_E_CTRL_INST_intermed_1 <= R.E.CTRL.INST;
		R_E_CTRL_INST_intermed_2 <= R_E_CTRL_INST_intermed_1;
		R_M_CTRL_INST_intermed_1 <= R.M.CTRL.INST;
		DE_INST_shadow_intermed_1 <= DE_INST_shadow;
		DE_INST_shadow_intermed_2 <= DE_INST_shadow_intermed_1;
		DE_INST_shadow_intermed_3 <= DE_INST_shadow_intermed_2;
		DE_INST_shadow_intermed_4 <= DE_INST_shadow_intermed_3;
		V_A_CTRL_INST_shadow_intermed_1 <= V_A_CTRL_INST_shadow;
		V_A_CTRL_INST_shadow_intermed_2 <= V_A_CTRL_INST_shadow_intermed_1;
		V_A_CTRL_INST_shadow_intermed_3 <= V_A_CTRL_INST_shadow_intermed_2;
		V_A_CTRL_INST_shadow_intermed_4 <= V_A_CTRL_INST_shadow_intermed_3;
		V_E_CTRL_INST_shadow_intermed_1 <= V_E_CTRL_INST_shadow;
		V_E_CTRL_INST_shadow_intermed_2 <= V_E_CTRL_INST_shadow_intermed_1;
		V_E_CTRL_INST_shadow_intermed_3 <= V_E_CTRL_INST_shadow_intermed_2;
		RIN_X_CTRL_INST_intermed_1 <= RIN.X.CTRL.INST;
		RIN_A_CTRL_INST_intermed_1 <= RIN.A.CTRL.INST;
		RIN_A_CTRL_INST_intermed_2 <= RIN_A_CTRL_INST_intermed_1;
		RIN_A_CTRL_INST_intermed_3 <= RIN_A_CTRL_INST_intermed_2;
		RIN_A_CTRL_INST_intermed_4 <= RIN_A_CTRL_INST_intermed_3;
		RIN_M_CTRL_INST_intermed_1 <= RIN.M.CTRL.INST;
		RIN_M_CTRL_INST_intermed_2 <= RIN_M_CTRL_INST_intermed_1;
		RIN_E_CTRL_INST_intermed_1 <= RIN.E.CTRL.INST;
		RIN_E_CTRL_INST_intermed_2 <= RIN_E_CTRL_INST_intermed_1;
		RIN_E_CTRL_INST_intermed_3 <= RIN_E_CTRL_INST_intermed_2;
		V_M_CTRL_INST_shadow_intermed_1 <= V_M_CTRL_INST_shadow;
		V_M_CTRL_INST_shadow_intermed_2 <= V_M_CTRL_INST_shadow_intermed_1;
		R_A_CTRL_INST_intermed_1 <= R.A.CTRL.INST;
		R_A_CTRL_INST_intermed_2 <= R_A_CTRL_INST_intermed_1;
		R_A_CTRL_INST_intermed_3 <= R_A_CTRL_INST_intermed_2;
		V_E_CTRL_CNT_shadow_intermed_1 <= V_E_CTRL_CNT_shadow;
		V_E_CTRL_CNT_shadow_intermed_2 <= V_E_CTRL_CNT_shadow_intermed_1;
		V_E_CTRL_CNT_shadow_intermed_3 <= V_E_CTRL_CNT_shadow_intermed_2;
		RIN_D_CNT_intermed_1 <= RIN.D.CNT;
		RIN_D_CNT_intermed_2 <= RIN_D_CNT_intermed_1;
		RIN_D_CNT_intermed_3 <= RIN_D_CNT_intermed_2;
		RIN_D_CNT_intermed_4 <= RIN_D_CNT_intermed_3;
		RIN_D_CNT_intermed_5 <= RIN_D_CNT_intermed_4;
		R_M_CTRL_CNT_intermed_1 <= R.M.CTRL.CNT;
		V_A_CTRL_CNT_shadow_intermed_1 <= V_A_CTRL_CNT_shadow;
		V_A_CTRL_CNT_shadow_intermed_2 <= V_A_CTRL_CNT_shadow_intermed_1;
		V_A_CTRL_CNT_shadow_intermed_3 <= V_A_CTRL_CNT_shadow_intermed_2;
		V_A_CTRL_CNT_shadow_intermed_4 <= V_A_CTRL_CNT_shadow_intermed_3;
		R_A_CTRL_CNT_intermed_1 <= R.A.CTRL.CNT;
		R_A_CTRL_CNT_intermed_2 <= R_A_CTRL_CNT_intermed_1;
		R_A_CTRL_CNT_intermed_3 <= R_A_CTRL_CNT_intermed_2;
		V_D_CNT_shadow_intermed_1 <= V_D_CNT_shadow;
		V_D_CNT_shadow_intermed_2 <= V_D_CNT_shadow_intermed_1;
		V_D_CNT_shadow_intermed_3 <= V_D_CNT_shadow_intermed_2;
		V_D_CNT_shadow_intermed_4 <= V_D_CNT_shadow_intermed_3;
		V_D_CNT_shadow_intermed_5 <= V_D_CNT_shadow_intermed_4;
		R_D_CNT_intermed_1 <= R.D.CNT;
		R_D_CNT_intermed_2 <= R_D_CNT_intermed_1;
		R_D_CNT_intermed_3 <= R_D_CNT_intermed_2;
		R_D_CNT_intermed_4 <= R_D_CNT_intermed_3;
		R_E_CTRL_CNT_intermed_1 <= R.E.CTRL.CNT;
		R_E_CTRL_CNT_intermed_2 <= R_E_CTRL_CNT_intermed_1;
		RIN_X_CTRL_CNT_intermed_1 <= RIN.X.CTRL.CNT;
		RIN_A_CTRL_CNT_intermed_1 <= RIN.A.CTRL.CNT;
		RIN_A_CTRL_CNT_intermed_2 <= RIN_A_CTRL_CNT_intermed_1;
		RIN_A_CTRL_CNT_intermed_3 <= RIN_A_CTRL_CNT_intermed_2;
		RIN_A_CTRL_CNT_intermed_4 <= RIN_A_CTRL_CNT_intermed_3;
		RIN_M_CTRL_CNT_intermed_1 <= RIN.M.CTRL.CNT;
		RIN_M_CTRL_CNT_intermed_2 <= RIN_M_CTRL_CNT_intermed_1;
		RIN_E_CTRL_CNT_intermed_1 <= RIN.E.CTRL.CNT;
		RIN_E_CTRL_CNT_intermed_2 <= RIN_E_CTRL_CNT_intermed_1;
		RIN_E_CTRL_CNT_intermed_3 <= RIN_E_CTRL_CNT_intermed_2;
		V_M_CTRL_CNT_shadow_intermed_1 <= V_M_CTRL_CNT_shadow;
		V_M_CTRL_CNT_shadow_intermed_2 <= V_M_CTRL_CNT_shadow_intermed_1;
		V_E_CTRL_PV_shadow_intermed_1 <= V_E_CTRL_PV_shadow;
		V_E_CTRL_PV_shadow_intermed_2 <= V_E_CTRL_PV_shadow_intermed_1;
		V_E_CTRL_PV_shadow_intermed_3 <= V_E_CTRL_PV_shadow_intermed_2;
		R_M_CTRL_PV_intermed_1 <= R.M.CTRL.PV;
		R_E_CTRL_PV_intermed_1 <= R.E.CTRL.PV;
		R_E_CTRL_PV_intermed_2 <= R_E_CTRL_PV_intermed_1;
		R_A_CTRL_PV_intermed_1 <= R.A.CTRL.PV;
		R_A_CTRL_PV_intermed_2 <= R_A_CTRL_PV_intermed_1;
		R_A_CTRL_PV_intermed_3 <= R_A_CTRL_PV_intermed_2;
		RIN_E_CTRL_PV_intermed_1 <= RIN.E.CTRL.PV;
		RIN_E_CTRL_PV_intermed_2 <= RIN_E_CTRL_PV_intermed_1;
		RIN_E_CTRL_PV_intermed_3 <= RIN_E_CTRL_PV_intermed_2;
		RIN_X_CTRL_PV_intermed_1 <= RIN.X.CTRL.PV;
		RIN_M_CTRL_PV_intermed_1 <= RIN.M.CTRL.PV;
		RIN_M_CTRL_PV_intermed_2 <= RIN_M_CTRL_PV_intermed_1;
		V_A_CTRL_PV_shadow_intermed_1 <= V_A_CTRL_PV_shadow;
		V_A_CTRL_PV_shadow_intermed_2 <= V_A_CTRL_PV_shadow_intermed_1;
		V_A_CTRL_PV_shadow_intermed_3 <= V_A_CTRL_PV_shadow_intermed_2;
		V_A_CTRL_PV_shadow_intermed_4 <= V_A_CTRL_PV_shadow_intermed_3;
		V_M_CTRL_PV_shadow_intermed_1 <= V_M_CTRL_PV_shadow;
		V_M_CTRL_PV_shadow_intermed_2 <= V_M_CTRL_PV_shadow_intermed_1;
		RIN_A_CTRL_PV_intermed_1 <= RIN.A.CTRL.PV;
		RIN_A_CTRL_PV_intermed_2 <= RIN_A_CTRL_PV_intermed_1;
		RIN_A_CTRL_PV_intermed_3 <= RIN_A_CTRL_PV_intermed_2;
		RIN_A_CTRL_PV_intermed_4 <= RIN_A_CTRL_PV_intermed_3;
		V_A_CTRL_INST19_shadow_intermed_1 <= V_A_CTRL_INST19_shadow;
		V_A_CTRL_INST19_shadow_intermed_2 <= V_A_CTRL_INST19_shadow_intermed_1;
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST( 19 );
		RIN_A_CTRL_INST19_intermed_2 <= RIN_A_CTRL_INST19_intermed_1;
		RIN_E_CTRL_INST19_intermed_1 <= RIN.E.CTRL.INST( 19 );
		DE_INST19_shadow_intermed_1 <= DE_INST19_shadow;
		DE_INST19_shadow_intermed_2 <= DE_INST19_shadow_intermed_1;
		R_A_CTRL_INST19_intermed_1 <= R.A.CTRL.INST( 19 );
		RIN_A_CTRL_INST20_intermed_1 <= RIN.A.CTRL.INST( 20 );
		RIN_A_CTRL_INST20_intermed_2 <= RIN_A_CTRL_INST20_intermed_1;
		V_A_CTRL_INST20_shadow_intermed_1 <= V_A_CTRL_INST20_shadow;
		V_A_CTRL_INST20_shadow_intermed_2 <= V_A_CTRL_INST20_shadow_intermed_1;
		RIN_E_CTRL_INST20_intermed_1 <= RIN.E.CTRL.INST( 20 );
		DE_INST20_shadow_intermed_1 <= DE_INST20_shadow;
		DE_INST20_shadow_intermed_2 <= DE_INST20_shadow_intermed_1;
		R_A_CTRL_INST20_intermed_1 <= R.A.CTRL.INST( 20 );
		R_A_CTRL_INST24_intermed_1 <= R.A.CTRL.INST( 24 );
		RIN_A_CTRL_INST24_intermed_1 <= RIN.A.CTRL.INST( 24 );
		RIN_A_CTRL_INST24_intermed_2 <= RIN_A_CTRL_INST24_intermed_1;
		RIN_E_CTRL_INST24_intermed_1 <= RIN.E.CTRL.INST( 24 );
		V_A_CTRL_INST24_shadow_intermed_1 <= V_A_CTRL_INST24_shadow;
		V_A_CTRL_INST24_shadow_intermed_2 <= V_A_CTRL_INST24_shadow_intermed_1;
		DE_INST24_shadow_intermed_1 <= DE_INST24_shadow;
		DE_INST24_shadow_intermed_2 <= DE_INST24_shadow_intermed_1;
		RIN_A_CTRL_INST19_intermed_1 <= RIN.A.CTRL.INST( 19 );
		DE_INST19_shadow_intermed_1 <= DE_INST19_shadow;
		V_X_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO4_shadow;
		V_X_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO4_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO4_shadow_intermed_3 <= V_X_CTRL_PC31DOWNTO4_shadow_intermed_2;
		IR_ADDR31DOWNTO4_intermed_1 <= IR.ADDR( 31 DOWNTO 4 );
		VIR_ADDR31DOWNTO4_shadow_intermed_1 <= VIR_ADDR31DOWNTO4_shadow;
		VIR_ADDR31DOWNTO4_shadow_intermed_2 <= VIR_ADDR31DOWNTO4_shadow_intermed_1;
		RIN_F_PC31DOWNTO4_intermed_1 <= RIN.F.PC( 31 DOWNTO 4 );
		RIN_A_CTRL_PC31DOWNTO4_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 4 );
		RIN_A_CTRL_PC31DOWNTO4_intermed_2 <= RIN_A_CTRL_PC31DOWNTO4_intermed_1;
		RIN_A_CTRL_PC31DOWNTO4_intermed_3 <= RIN_A_CTRL_PC31DOWNTO4_intermed_2;
		RIN_A_CTRL_PC31DOWNTO4_intermed_4 <= RIN_A_CTRL_PC31DOWNTO4_intermed_3;
		RIN_A_CTRL_PC31DOWNTO4_intermed_5 <= RIN_A_CTRL_PC31DOWNTO4_intermed_4;
		RIN_A_CTRL_PC31DOWNTO4_intermed_6 <= RIN_A_CTRL_PC31DOWNTO4_intermed_5;
		R_A_CTRL_PC31DOWNTO4_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 4 );
		R_A_CTRL_PC31DOWNTO4_intermed_2 <= R_A_CTRL_PC31DOWNTO4_intermed_1;
		R_A_CTRL_PC31DOWNTO4_intermed_3 <= R_A_CTRL_PC31DOWNTO4_intermed_2;
		R_A_CTRL_PC31DOWNTO4_intermed_4 <= R_A_CTRL_PC31DOWNTO4_intermed_3;
		R_A_CTRL_PC31DOWNTO4_intermed_5 <= R_A_CTRL_PC31DOWNTO4_intermed_4;
		R_D_PC31DOWNTO4_intermed_1 <= R.D.PC( 31 DOWNTO 4 );
		R_D_PC31DOWNTO4_intermed_2 <= R_D_PC31DOWNTO4_intermed_1;
		R_D_PC31DOWNTO4_intermed_3 <= R_D_PC31DOWNTO4_intermed_2;
		R_D_PC31DOWNTO4_intermed_4 <= R_D_PC31DOWNTO4_intermed_3;
		R_D_PC31DOWNTO4_intermed_5 <= R_D_PC31DOWNTO4_intermed_4;
		R_D_PC31DOWNTO4_intermed_6 <= R_D_PC31DOWNTO4_intermed_5;
		RIN_X_CTRL_PC31DOWNTO4_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 4 );
		RIN_X_CTRL_PC31DOWNTO4_intermed_2 <= RIN_X_CTRL_PC31DOWNTO4_intermed_1;
		RIN_X_CTRL_PC31DOWNTO4_intermed_3 <= RIN_X_CTRL_PC31DOWNTO4_intermed_2;
		EX_ADD_RES32DOWNTO332DOWNTO5_shadow_intermed_1 <= EX_ADD_RES32DOWNTO332DOWNTO5_shadow;
		V_D_PC31DOWNTO4_shadow_intermed_1 <= V_D_PC31DOWNTO4_shadow;
		V_D_PC31DOWNTO4_shadow_intermed_2 <= V_D_PC31DOWNTO4_shadow_intermed_1;
		V_D_PC31DOWNTO4_shadow_intermed_3 <= V_D_PC31DOWNTO4_shadow_intermed_2;
		V_D_PC31DOWNTO4_shadow_intermed_4 <= V_D_PC31DOWNTO4_shadow_intermed_3;
		V_D_PC31DOWNTO4_shadow_intermed_5 <= V_D_PC31DOWNTO4_shadow_intermed_4;
		V_D_PC31DOWNTO4_shadow_intermed_6 <= V_D_PC31DOWNTO4_shadow_intermed_5;
		V_D_PC31DOWNTO4_shadow_intermed_7 <= V_D_PC31DOWNTO4_shadow_intermed_6;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO4_shadow;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO4_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO4_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO4_shadow_intermed_3;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_5 <= V_E_CTRL_PC31DOWNTO4_shadow_intermed_4;
		RIN_M_CTRL_PC31DOWNTO4_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 4 );
		RIN_M_CTRL_PC31DOWNTO4_intermed_2 <= RIN_M_CTRL_PC31DOWNTO4_intermed_1;
		RIN_M_CTRL_PC31DOWNTO4_intermed_3 <= RIN_M_CTRL_PC31DOWNTO4_intermed_2;
		RIN_M_CTRL_PC31DOWNTO4_intermed_4 <= RIN_M_CTRL_PC31DOWNTO4_intermed_3;
		R_X_CTRL_PC31DOWNTO4_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 4 );
		R_X_CTRL_PC31DOWNTO4_intermed_2 <= R_X_CTRL_PC31DOWNTO4_intermed_1;
		IRIN_ADDR31DOWNTO4_intermed_1 <= IRIN.ADDR( 31 DOWNTO 4 );
		IRIN_ADDR31DOWNTO4_intermed_2 <= IRIN_ADDR31DOWNTO4_intermed_1;
		V_M_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO4_shadow;
		V_M_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO4_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO4_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO4_shadow_intermed_2;
		V_M_CTRL_PC31DOWNTO4_shadow_intermed_4 <= V_M_CTRL_PC31DOWNTO4_shadow_intermed_3;
		R_M_CTRL_PC31DOWNTO4_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 4 );
		R_M_CTRL_PC31DOWNTO4_intermed_2 <= R_M_CTRL_PC31DOWNTO4_intermed_1;
		R_M_CTRL_PC31DOWNTO4_intermed_3 <= R_M_CTRL_PC31DOWNTO4_intermed_2;
		XC_TRAP_ADDRESS31DOWNTO4_shadow_intermed_1 <= XC_TRAP_ADDRESS31DOWNTO4_shadow;
		RIN_D_PC31DOWNTO4_intermed_1 <= RIN.D.PC( 31 DOWNTO 4 );
		RIN_D_PC31DOWNTO4_intermed_2 <= RIN_D_PC31DOWNTO4_intermed_1;
		RIN_D_PC31DOWNTO4_intermed_3 <= RIN_D_PC31DOWNTO4_intermed_2;
		RIN_D_PC31DOWNTO4_intermed_4 <= RIN_D_PC31DOWNTO4_intermed_3;
		RIN_D_PC31DOWNTO4_intermed_5 <= RIN_D_PC31DOWNTO4_intermed_4;
		RIN_D_PC31DOWNTO4_intermed_6 <= RIN_D_PC31DOWNTO4_intermed_5;
		RIN_D_PC31DOWNTO4_intermed_7 <= RIN_D_PC31DOWNTO4_intermed_6;
		RIN_E_CTRL_PC31DOWNTO4_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 4 );
		RIN_E_CTRL_PC31DOWNTO4_intermed_2 <= RIN_E_CTRL_PC31DOWNTO4_intermed_1;
		RIN_E_CTRL_PC31DOWNTO4_intermed_3 <= RIN_E_CTRL_PC31DOWNTO4_intermed_2;
		RIN_E_CTRL_PC31DOWNTO4_intermed_4 <= RIN_E_CTRL_PC31DOWNTO4_intermed_3;
		RIN_E_CTRL_PC31DOWNTO4_intermed_5 <= RIN_E_CTRL_PC31DOWNTO4_intermed_4;
		EX_JUMP_ADDRESS31DOWNTO4_shadow_intermed_1 <= EX_JUMP_ADDRESS31DOWNTO4_shadow;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO4_shadow;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_4;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_6 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_5;
		R_E_CTRL_PC31DOWNTO4_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 4 );
		R_E_CTRL_PC31DOWNTO4_intermed_2 <= R_E_CTRL_PC31DOWNTO4_intermed_1;
		R_E_CTRL_PC31DOWNTO4_intermed_3 <= R_E_CTRL_PC31DOWNTO4_intermed_2;
		R_E_CTRL_PC31DOWNTO4_intermed_4 <= R_E_CTRL_PC31DOWNTO4_intermed_3;
		V_X_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO4_shadow;
		V_X_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO4_shadow_intermed_1;
		RIN_A_CTRL_PC31DOWNTO4_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 4 );
		RIN_A_CTRL_PC31DOWNTO4_intermed_2 <= RIN_A_CTRL_PC31DOWNTO4_intermed_1;
		RIN_A_CTRL_PC31DOWNTO4_intermed_3 <= RIN_A_CTRL_PC31DOWNTO4_intermed_2;
		RIN_A_CTRL_PC31DOWNTO4_intermed_4 <= RIN_A_CTRL_PC31DOWNTO4_intermed_3;
		RIN_A_CTRL_PC31DOWNTO4_intermed_5 <= RIN_A_CTRL_PC31DOWNTO4_intermed_4;
		R_A_CTRL_PC31DOWNTO4_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 4 );
		R_A_CTRL_PC31DOWNTO4_intermed_2 <= R_A_CTRL_PC31DOWNTO4_intermed_1;
		R_A_CTRL_PC31DOWNTO4_intermed_3 <= R_A_CTRL_PC31DOWNTO4_intermed_2;
		R_A_CTRL_PC31DOWNTO4_intermed_4 <= R_A_CTRL_PC31DOWNTO4_intermed_3;
		R_D_PC31DOWNTO4_intermed_1 <= R.D.PC( 31 DOWNTO 4 );
		R_D_PC31DOWNTO4_intermed_2 <= R_D_PC31DOWNTO4_intermed_1;
		R_D_PC31DOWNTO4_intermed_3 <= R_D_PC31DOWNTO4_intermed_2;
		R_D_PC31DOWNTO4_intermed_4 <= R_D_PC31DOWNTO4_intermed_3;
		R_D_PC31DOWNTO4_intermed_5 <= R_D_PC31DOWNTO4_intermed_4;
		RIN_X_CTRL_PC31DOWNTO4_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 4 );
		RIN_X_CTRL_PC31DOWNTO4_intermed_2 <= RIN_X_CTRL_PC31DOWNTO4_intermed_1;
		V_D_PC31DOWNTO4_shadow_intermed_1 <= V_D_PC31DOWNTO4_shadow;
		V_D_PC31DOWNTO4_shadow_intermed_2 <= V_D_PC31DOWNTO4_shadow_intermed_1;
		V_D_PC31DOWNTO4_shadow_intermed_3 <= V_D_PC31DOWNTO4_shadow_intermed_2;
		V_D_PC31DOWNTO4_shadow_intermed_4 <= V_D_PC31DOWNTO4_shadow_intermed_3;
		V_D_PC31DOWNTO4_shadow_intermed_5 <= V_D_PC31DOWNTO4_shadow_intermed_4;
		V_D_PC31DOWNTO4_shadow_intermed_6 <= V_D_PC31DOWNTO4_shadow_intermed_5;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO4_shadow;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO4_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO4_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO4_shadow_intermed_3;
		RIN_M_CTRL_PC31DOWNTO4_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 4 );
		RIN_M_CTRL_PC31DOWNTO4_intermed_2 <= RIN_M_CTRL_PC31DOWNTO4_intermed_1;
		RIN_M_CTRL_PC31DOWNTO4_intermed_3 <= RIN_M_CTRL_PC31DOWNTO4_intermed_2;
		R_X_CTRL_PC31DOWNTO4_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 4 );
		IRIN_ADDR31DOWNTO4_intermed_1 <= IRIN.ADDR( 31 DOWNTO 4 );
		V_M_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO4_shadow;
		V_M_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO4_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO4_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO4_shadow_intermed_2;
		R_M_CTRL_PC31DOWNTO4_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 4 );
		R_M_CTRL_PC31DOWNTO4_intermed_2 <= R_M_CTRL_PC31DOWNTO4_intermed_1;
		RIN_D_PC31DOWNTO4_intermed_1 <= RIN.D.PC( 31 DOWNTO 4 );
		RIN_D_PC31DOWNTO4_intermed_2 <= RIN_D_PC31DOWNTO4_intermed_1;
		RIN_D_PC31DOWNTO4_intermed_3 <= RIN_D_PC31DOWNTO4_intermed_2;
		RIN_D_PC31DOWNTO4_intermed_4 <= RIN_D_PC31DOWNTO4_intermed_3;
		RIN_D_PC31DOWNTO4_intermed_5 <= RIN_D_PC31DOWNTO4_intermed_4;
		RIN_D_PC31DOWNTO4_intermed_6 <= RIN_D_PC31DOWNTO4_intermed_5;
		RIN_E_CTRL_PC31DOWNTO4_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 4 );
		RIN_E_CTRL_PC31DOWNTO4_intermed_2 <= RIN_E_CTRL_PC31DOWNTO4_intermed_1;
		RIN_E_CTRL_PC31DOWNTO4_intermed_3 <= RIN_E_CTRL_PC31DOWNTO4_intermed_2;
		RIN_E_CTRL_PC31DOWNTO4_intermed_4 <= RIN_E_CTRL_PC31DOWNTO4_intermed_3;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO4_shadow;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_4;
		R_E_CTRL_PC31DOWNTO4_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 4 );
		R_E_CTRL_PC31DOWNTO4_intermed_2 <= R_E_CTRL_PC31DOWNTO4_intermed_1;
		R_E_CTRL_PC31DOWNTO4_intermed_3 <= R_E_CTRL_PC31DOWNTO4_intermed_2;
		R_D_PC3DOWNTO2_intermed_1 <= R.D.PC( 3 DOWNTO 2 );
		R_D_PC3DOWNTO2_intermed_2 <= R_D_PC3DOWNTO2_intermed_1;
		R_D_PC3DOWNTO2_intermed_3 <= R_D_PC3DOWNTO2_intermed_2;
		R_D_PC3DOWNTO2_intermed_4 <= R_D_PC3DOWNTO2_intermed_3;
		R_D_PC3DOWNTO2_intermed_5 <= R_D_PC3DOWNTO2_intermed_4;
		R_D_PC3DOWNTO2_intermed_6 <= R_D_PC3DOWNTO2_intermed_5;
		V_D_PC3DOWNTO2_shadow_intermed_1 <= V_D_PC3DOWNTO2_shadow;
		V_D_PC3DOWNTO2_shadow_intermed_2 <= V_D_PC3DOWNTO2_shadow_intermed_1;
		V_D_PC3DOWNTO2_shadow_intermed_3 <= V_D_PC3DOWNTO2_shadow_intermed_2;
		V_D_PC3DOWNTO2_shadow_intermed_4 <= V_D_PC3DOWNTO2_shadow_intermed_3;
		V_D_PC3DOWNTO2_shadow_intermed_5 <= V_D_PC3DOWNTO2_shadow_intermed_4;
		V_D_PC3DOWNTO2_shadow_intermed_6 <= V_D_PC3DOWNTO2_shadow_intermed_5;
		V_D_PC3DOWNTO2_shadow_intermed_7 <= V_D_PC3DOWNTO2_shadow_intermed_6;
		VIR_ADDR3DOWNTO2_shadow_intermed_1 <= VIR_ADDR3DOWNTO2_shadow;
		VIR_ADDR3DOWNTO2_shadow_intermed_2 <= VIR_ADDR3DOWNTO2_shadow_intermed_1;
		RIN_D_PC3DOWNTO2_intermed_1 <= RIN.D.PC( 3 DOWNTO 2 );
		RIN_D_PC3DOWNTO2_intermed_2 <= RIN_D_PC3DOWNTO2_intermed_1;
		RIN_D_PC3DOWNTO2_intermed_3 <= RIN_D_PC3DOWNTO2_intermed_2;
		RIN_D_PC3DOWNTO2_intermed_4 <= RIN_D_PC3DOWNTO2_intermed_3;
		RIN_D_PC3DOWNTO2_intermed_5 <= RIN_D_PC3DOWNTO2_intermed_4;
		RIN_D_PC3DOWNTO2_intermed_6 <= RIN_D_PC3DOWNTO2_intermed_5;
		RIN_D_PC3DOWNTO2_intermed_7 <= RIN_D_PC3DOWNTO2_intermed_6;
		R_M_CTRL_PC3DOWNTO2_intermed_1 <= R.M.CTRL.PC( 3 DOWNTO 2 );
		R_M_CTRL_PC3DOWNTO2_intermed_2 <= R_M_CTRL_PC3DOWNTO2_intermed_1;
		R_M_CTRL_PC3DOWNTO2_intermed_3 <= R_M_CTRL_PC3DOWNTO2_intermed_2;
		R_E_CTRL_PC3DOWNTO2_intermed_1 <= R.E.CTRL.PC( 3 DOWNTO 2 );
		R_E_CTRL_PC3DOWNTO2_intermed_2 <= R_E_CTRL_PC3DOWNTO2_intermed_1;
		R_E_CTRL_PC3DOWNTO2_intermed_3 <= R_E_CTRL_PC3DOWNTO2_intermed_2;
		R_E_CTRL_PC3DOWNTO2_intermed_4 <= R_E_CTRL_PC3DOWNTO2_intermed_3;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC3DOWNTO2_shadow;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC3DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC3DOWNTO2_shadow_intermed_2;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_4 <= V_E_CTRL_PC3DOWNTO2_shadow_intermed_3;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_5 <= V_E_CTRL_PC3DOWNTO2_shadow_intermed_4;
		RIN_X_CTRL_PC3DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 3 DOWNTO 2 );
		RIN_X_CTRL_PC3DOWNTO2_intermed_2 <= RIN_X_CTRL_PC3DOWNTO2_intermed_1;
		RIN_X_CTRL_PC3DOWNTO2_intermed_3 <= RIN_X_CTRL_PC3DOWNTO2_intermed_2;
		R_A_CTRL_PC3DOWNTO2_intermed_1 <= R.A.CTRL.PC( 3 DOWNTO 2 );
		R_A_CTRL_PC3DOWNTO2_intermed_2 <= R_A_CTRL_PC3DOWNTO2_intermed_1;
		R_A_CTRL_PC3DOWNTO2_intermed_3 <= R_A_CTRL_PC3DOWNTO2_intermed_2;
		R_A_CTRL_PC3DOWNTO2_intermed_4 <= R_A_CTRL_PC3DOWNTO2_intermed_3;
		R_A_CTRL_PC3DOWNTO2_intermed_5 <= R_A_CTRL_PC3DOWNTO2_intermed_4;
		V_X_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC3DOWNTO2_shadow;
		V_X_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_X_CTRL_PC3DOWNTO2_shadow_intermed_1;
		V_X_CTRL_PC3DOWNTO2_shadow_intermed_3 <= V_X_CTRL_PC3DOWNTO2_shadow_intermed_2;
		RIN_M_CTRL_PC3DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 3 DOWNTO 2 );
		RIN_M_CTRL_PC3DOWNTO2_intermed_2 <= RIN_M_CTRL_PC3DOWNTO2_intermed_1;
		RIN_M_CTRL_PC3DOWNTO2_intermed_3 <= RIN_M_CTRL_PC3DOWNTO2_intermed_2;
		RIN_M_CTRL_PC3DOWNTO2_intermed_4 <= RIN_M_CTRL_PC3DOWNTO2_intermed_3;
		IRIN_ADDR3DOWNTO2_intermed_1 <= IRIN.ADDR( 3 DOWNTO 2 );
		IRIN_ADDR3DOWNTO2_intermed_2 <= IRIN_ADDR3DOWNTO2_intermed_1;
		EX_JUMP_ADDRESS3DOWNTO2_shadow_intermed_1 <= EX_JUMP_ADDRESS3DOWNTO2_shadow;
		EX_ADD_RES32DOWNTO34DOWNTO3_shadow_intermed_1 <= EX_ADD_RES32DOWNTO34DOWNTO3_shadow;
		RIN_A_CTRL_PC3DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 3 DOWNTO 2 );
		RIN_A_CTRL_PC3DOWNTO2_intermed_2 <= RIN_A_CTRL_PC3DOWNTO2_intermed_1;
		RIN_A_CTRL_PC3DOWNTO2_intermed_3 <= RIN_A_CTRL_PC3DOWNTO2_intermed_2;
		RIN_A_CTRL_PC3DOWNTO2_intermed_4 <= RIN_A_CTRL_PC3DOWNTO2_intermed_3;
		RIN_A_CTRL_PC3DOWNTO2_intermed_5 <= RIN_A_CTRL_PC3DOWNTO2_intermed_4;
		RIN_A_CTRL_PC3DOWNTO2_intermed_6 <= RIN_A_CTRL_PC3DOWNTO2_intermed_5;
		XC_TRAP_ADDRESS3DOWNTO2_shadow_intermed_1 <= XC_TRAP_ADDRESS3DOWNTO2_shadow;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC3DOWNTO2_shadow;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_3;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_5 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_4;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_6 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_5;
		IR_ADDR3DOWNTO2_intermed_1 <= IR.ADDR( 3 DOWNTO 2 );
		V_M_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC3DOWNTO2_shadow;
		V_M_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC3DOWNTO2_shadow_intermed_1;
		V_M_CTRL_PC3DOWNTO2_shadow_intermed_3 <= V_M_CTRL_PC3DOWNTO2_shadow_intermed_2;
		V_M_CTRL_PC3DOWNTO2_shadow_intermed_4 <= V_M_CTRL_PC3DOWNTO2_shadow_intermed_3;
		R_X_CTRL_PC3DOWNTO2_intermed_1 <= R.X.CTRL.PC( 3 DOWNTO 2 );
		R_X_CTRL_PC3DOWNTO2_intermed_2 <= R_X_CTRL_PC3DOWNTO2_intermed_1;
		RIN_E_CTRL_PC3DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 3 DOWNTO 2 );
		RIN_E_CTRL_PC3DOWNTO2_intermed_2 <= RIN_E_CTRL_PC3DOWNTO2_intermed_1;
		RIN_E_CTRL_PC3DOWNTO2_intermed_3 <= RIN_E_CTRL_PC3DOWNTO2_intermed_2;
		RIN_E_CTRL_PC3DOWNTO2_intermed_4 <= RIN_E_CTRL_PC3DOWNTO2_intermed_3;
		RIN_E_CTRL_PC3DOWNTO2_intermed_5 <= RIN_E_CTRL_PC3DOWNTO2_intermed_4;
		RIN_F_PC3DOWNTO2_intermed_1 <= RIN.F.PC( 3 DOWNTO 2 );
		R_D_PC3DOWNTO2_intermed_1 <= R.D.PC( 3 DOWNTO 2 );
		R_D_PC3DOWNTO2_intermed_2 <= R_D_PC3DOWNTO2_intermed_1;
		R_D_PC3DOWNTO2_intermed_3 <= R_D_PC3DOWNTO2_intermed_2;
		R_D_PC3DOWNTO2_intermed_4 <= R_D_PC3DOWNTO2_intermed_3;
		R_D_PC3DOWNTO2_intermed_5 <= R_D_PC3DOWNTO2_intermed_4;
		V_D_PC3DOWNTO2_shadow_intermed_1 <= V_D_PC3DOWNTO2_shadow;
		V_D_PC3DOWNTO2_shadow_intermed_2 <= V_D_PC3DOWNTO2_shadow_intermed_1;
		V_D_PC3DOWNTO2_shadow_intermed_3 <= V_D_PC3DOWNTO2_shadow_intermed_2;
		V_D_PC3DOWNTO2_shadow_intermed_4 <= V_D_PC3DOWNTO2_shadow_intermed_3;
		V_D_PC3DOWNTO2_shadow_intermed_5 <= V_D_PC3DOWNTO2_shadow_intermed_4;
		V_D_PC3DOWNTO2_shadow_intermed_6 <= V_D_PC3DOWNTO2_shadow_intermed_5;
		RIN_D_PC3DOWNTO2_intermed_1 <= RIN.D.PC( 3 DOWNTO 2 );
		RIN_D_PC3DOWNTO2_intermed_2 <= RIN_D_PC3DOWNTO2_intermed_1;
		RIN_D_PC3DOWNTO2_intermed_3 <= RIN_D_PC3DOWNTO2_intermed_2;
		RIN_D_PC3DOWNTO2_intermed_4 <= RIN_D_PC3DOWNTO2_intermed_3;
		RIN_D_PC3DOWNTO2_intermed_5 <= RIN_D_PC3DOWNTO2_intermed_4;
		RIN_D_PC3DOWNTO2_intermed_6 <= RIN_D_PC3DOWNTO2_intermed_5;
		R_M_CTRL_PC3DOWNTO2_intermed_1 <= R.M.CTRL.PC( 3 DOWNTO 2 );
		R_M_CTRL_PC3DOWNTO2_intermed_2 <= R_M_CTRL_PC3DOWNTO2_intermed_1;
		R_E_CTRL_PC3DOWNTO2_intermed_1 <= R.E.CTRL.PC( 3 DOWNTO 2 );
		R_E_CTRL_PC3DOWNTO2_intermed_2 <= R_E_CTRL_PC3DOWNTO2_intermed_1;
		R_E_CTRL_PC3DOWNTO2_intermed_3 <= R_E_CTRL_PC3DOWNTO2_intermed_2;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC3DOWNTO2_shadow;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC3DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC3DOWNTO2_shadow_intermed_2;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_4 <= V_E_CTRL_PC3DOWNTO2_shadow_intermed_3;
		RIN_X_CTRL_PC3DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 3 DOWNTO 2 );
		RIN_X_CTRL_PC3DOWNTO2_intermed_2 <= RIN_X_CTRL_PC3DOWNTO2_intermed_1;
		R_A_CTRL_PC3DOWNTO2_intermed_1 <= R.A.CTRL.PC( 3 DOWNTO 2 );
		R_A_CTRL_PC3DOWNTO2_intermed_2 <= R_A_CTRL_PC3DOWNTO2_intermed_1;
		R_A_CTRL_PC3DOWNTO2_intermed_3 <= R_A_CTRL_PC3DOWNTO2_intermed_2;
		R_A_CTRL_PC3DOWNTO2_intermed_4 <= R_A_CTRL_PC3DOWNTO2_intermed_3;
		V_X_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC3DOWNTO2_shadow;
		V_X_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_X_CTRL_PC3DOWNTO2_shadow_intermed_1;
		RIN_M_CTRL_PC3DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 3 DOWNTO 2 );
		RIN_M_CTRL_PC3DOWNTO2_intermed_2 <= RIN_M_CTRL_PC3DOWNTO2_intermed_1;
		RIN_M_CTRL_PC3DOWNTO2_intermed_3 <= RIN_M_CTRL_PC3DOWNTO2_intermed_2;
		IRIN_ADDR3DOWNTO2_intermed_1 <= IRIN.ADDR( 3 DOWNTO 2 );
		RIN_A_CTRL_PC3DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 3 DOWNTO 2 );
		RIN_A_CTRL_PC3DOWNTO2_intermed_2 <= RIN_A_CTRL_PC3DOWNTO2_intermed_1;
		RIN_A_CTRL_PC3DOWNTO2_intermed_3 <= RIN_A_CTRL_PC3DOWNTO2_intermed_2;
		RIN_A_CTRL_PC3DOWNTO2_intermed_4 <= RIN_A_CTRL_PC3DOWNTO2_intermed_3;
		RIN_A_CTRL_PC3DOWNTO2_intermed_5 <= RIN_A_CTRL_PC3DOWNTO2_intermed_4;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC3DOWNTO2_shadow;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_3;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_5 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_4;
		V_M_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC3DOWNTO2_shadow;
		V_M_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC3DOWNTO2_shadow_intermed_1;
		V_M_CTRL_PC3DOWNTO2_shadow_intermed_3 <= V_M_CTRL_PC3DOWNTO2_shadow_intermed_2;
		R_X_CTRL_PC3DOWNTO2_intermed_1 <= R.X.CTRL.PC( 3 DOWNTO 2 );
		RIN_E_CTRL_PC3DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 3 DOWNTO 2 );
		RIN_E_CTRL_PC3DOWNTO2_intermed_2 <= RIN_E_CTRL_PC3DOWNTO2_intermed_1;
		RIN_E_CTRL_PC3DOWNTO2_intermed_3 <= RIN_E_CTRL_PC3DOWNTO2_intermed_2;
		RIN_E_CTRL_PC3DOWNTO2_intermed_4 <= RIN_E_CTRL_PC3DOWNTO2_intermed_3;
		RIN_E_CTRL_RD6DOWNTO0_intermed_1 <= RIN.E.CTRL.RD( 6 DOWNTO 0 );
		RIN_E_CTRL_RD6DOWNTO0_intermed_2 <= RIN_E_CTRL_RD6DOWNTO0_intermed_1;
		RIN_E_CTRL_RD6DOWNTO0_intermed_3 <= RIN_E_CTRL_RD6DOWNTO0_intermed_2;
		RIN_M_CTRL_RD6DOWNTO0_intermed_1 <= RIN.M.CTRL.RD( 6 DOWNTO 0 );
		RIN_M_CTRL_RD6DOWNTO0_intermed_2 <= RIN_M_CTRL_RD6DOWNTO0_intermed_1;
		RIN_X_CTRL_RD6DOWNTO0_intermed_1 <= RIN.X.CTRL.RD( 6 DOWNTO 0 );
		V_M_CTRL_RD6DOWNTO0_shadow_intermed_1 <= V_M_CTRL_RD6DOWNTO0_shadow;
		V_M_CTRL_RD6DOWNTO0_shadow_intermed_2 <= V_M_CTRL_RD6DOWNTO0_shadow_intermed_1;
		R_E_CTRL_RD6DOWNTO0_intermed_1 <= R.E.CTRL.RD( 6 DOWNTO 0 );
		R_E_CTRL_RD6DOWNTO0_intermed_2 <= R_E_CTRL_RD6DOWNTO0_intermed_1;
		V_E_CTRL_RD6DOWNTO0_shadow_intermed_1 <= V_E_CTRL_RD6DOWNTO0_shadow;
		V_E_CTRL_RD6DOWNTO0_shadow_intermed_2 <= V_E_CTRL_RD6DOWNTO0_shadow_intermed_1;
		V_E_CTRL_RD6DOWNTO0_shadow_intermed_3 <= V_E_CTRL_RD6DOWNTO0_shadow_intermed_2;
		V_A_CTRL_RD6DOWNTO0_shadow_intermed_1 <= V_A_CTRL_RD6DOWNTO0_shadow;
		V_A_CTRL_RD6DOWNTO0_shadow_intermed_2 <= V_A_CTRL_RD6DOWNTO0_shadow_intermed_1;
		V_A_CTRL_RD6DOWNTO0_shadow_intermed_3 <= V_A_CTRL_RD6DOWNTO0_shadow_intermed_2;
		V_A_CTRL_RD6DOWNTO0_shadow_intermed_4 <= V_A_CTRL_RD6DOWNTO0_shadow_intermed_3;
		R_A_CTRL_RD6DOWNTO0_intermed_1 <= R.A.CTRL.RD( 6 DOWNTO 0 );
		R_A_CTRL_RD6DOWNTO0_intermed_2 <= R_A_CTRL_RD6DOWNTO0_intermed_1;
		R_A_CTRL_RD6DOWNTO0_intermed_3 <= R_A_CTRL_RD6DOWNTO0_intermed_2;
		RIN_A_CTRL_RD6DOWNTO0_intermed_1 <= RIN.A.CTRL.RD( 6 DOWNTO 0 );
		RIN_A_CTRL_RD6DOWNTO0_intermed_2 <= RIN_A_CTRL_RD6DOWNTO0_intermed_1;
		RIN_A_CTRL_RD6DOWNTO0_intermed_3 <= RIN_A_CTRL_RD6DOWNTO0_intermed_2;
		RIN_A_CTRL_RD6DOWNTO0_intermed_4 <= RIN_A_CTRL_RD6DOWNTO0_intermed_3;
		R_M_CTRL_RD6DOWNTO0_intermed_1 <= R.M.CTRL.RD( 6 DOWNTO 0 );
		V_E_CTRL_TT_shadow_intermed_1 <= V_E_CTRL_TT_shadow;
		V_E_CTRL_TT_shadow_intermed_2 <= V_E_CTRL_TT_shadow_intermed_1;
		RIN_A_CTRL_TT_intermed_1 <= RIN.A.CTRL.TT;
		RIN_A_CTRL_TT_intermed_2 <= RIN_A_CTRL_TT_intermed_1;
		RIN_A_CTRL_TT_intermed_3 <= RIN_A_CTRL_TT_intermed_2;
		R_A_CTRL_TT_intermed_1 <= R.A.CTRL.TT;
		R_A_CTRL_TT_intermed_2 <= R_A_CTRL_TT_intermed_1;
		R_E_CTRL_TT_intermed_1 <= R.E.CTRL.TT;
		RIN_M_CTRL_TT_intermed_1 <= RIN.M.CTRL.TT;
		RIN_E_CTRL_TT_intermed_1 <= RIN.E.CTRL.TT;
		RIN_E_CTRL_TT_intermed_2 <= RIN_E_CTRL_TT_intermed_1;
		V_A_CTRL_TT_shadow_intermed_1 <= V_A_CTRL_TT_shadow;
		V_A_CTRL_TT_shadow_intermed_2 <= V_A_CTRL_TT_shadow_intermed_1;
		V_A_CTRL_TT_shadow_intermed_3 <= V_A_CTRL_TT_shadow_intermed_2;
		R_A_CTRL_LD_intermed_1 <= R.A.CTRL.LD;
		RIN_A_CTRL_LD_intermed_1 <= RIN.A.CTRL.LD;
		RIN_A_CTRL_LD_intermed_2 <= RIN_A_CTRL_LD_intermed_1;
		RIN_E_CTRL_LD_intermed_1 <= RIN.E.CTRL.LD;
		V_A_CTRL_LD_shadow_intermed_1 <= V_A_CTRL_LD_shadow;
		V_A_CTRL_LD_shadow_intermed_2 <= V_A_CTRL_LD_shadow_intermed_1;
		R_M_CTRL_PC31DOWNTO12_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 12 );
		R_M_CTRL_PC31DOWNTO12_intermed_2 <= R_M_CTRL_PC31DOWNTO12_intermed_1;
		R_M_CTRL_PC31DOWNTO12_intermed_3 <= R_M_CTRL_PC31DOWNTO12_intermed_2;
		V_D_PC31DOWNTO12_shadow_intermed_1 <= V_D_PC31DOWNTO12_shadow;
		V_D_PC31DOWNTO12_shadow_intermed_2 <= V_D_PC31DOWNTO12_shadow_intermed_1;
		V_D_PC31DOWNTO12_shadow_intermed_3 <= V_D_PC31DOWNTO12_shadow_intermed_2;
		V_D_PC31DOWNTO12_shadow_intermed_4 <= V_D_PC31DOWNTO12_shadow_intermed_3;
		V_D_PC31DOWNTO12_shadow_intermed_5 <= V_D_PC31DOWNTO12_shadow_intermed_4;
		V_D_PC31DOWNTO12_shadow_intermed_6 <= V_D_PC31DOWNTO12_shadow_intermed_5;
		V_D_PC31DOWNTO12_shadow_intermed_7 <= V_D_PC31DOWNTO12_shadow_intermed_6;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO12_shadow;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_4;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_6 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_5;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO12_shadow;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_3;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_5 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_4;
		EX_ADD_RES32DOWNTO330DOWNTO11_shadow_intermed_1 <= EX_ADD_RES32DOWNTO330DOWNTO11_shadow;
		RIN_F_PC31DOWNTO12_intermed_1 <= RIN.F.PC( 31 DOWNTO 12 );
		R_A_CTRL_PC31DOWNTO12_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 12 );
		R_A_CTRL_PC31DOWNTO12_intermed_2 <= R_A_CTRL_PC31DOWNTO12_intermed_1;
		R_A_CTRL_PC31DOWNTO12_intermed_3 <= R_A_CTRL_PC31DOWNTO12_intermed_2;
		R_A_CTRL_PC31DOWNTO12_intermed_4 <= R_A_CTRL_PC31DOWNTO12_intermed_3;
		R_A_CTRL_PC31DOWNTO12_intermed_5 <= R_A_CTRL_PC31DOWNTO12_intermed_4;
		R_E_CTRL_PC31DOWNTO12_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 12 );
		R_E_CTRL_PC31DOWNTO12_intermed_2 <= R_E_CTRL_PC31DOWNTO12_intermed_1;
		R_E_CTRL_PC31DOWNTO12_intermed_3 <= R_E_CTRL_PC31DOWNTO12_intermed_2;
		R_E_CTRL_PC31DOWNTO12_intermed_4 <= R_E_CTRL_PC31DOWNTO12_intermed_3;
		EX_JUMP_ADDRESS31DOWNTO12_shadow_intermed_1 <= EX_JUMP_ADDRESS31DOWNTO12_shadow;
		RIN_A_CTRL_PC31DOWNTO12_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 12 );
		RIN_A_CTRL_PC31DOWNTO12_intermed_2 <= RIN_A_CTRL_PC31DOWNTO12_intermed_1;
		RIN_A_CTRL_PC31DOWNTO12_intermed_3 <= RIN_A_CTRL_PC31DOWNTO12_intermed_2;
		RIN_A_CTRL_PC31DOWNTO12_intermed_4 <= RIN_A_CTRL_PC31DOWNTO12_intermed_3;
		RIN_A_CTRL_PC31DOWNTO12_intermed_5 <= RIN_A_CTRL_PC31DOWNTO12_intermed_4;
		RIN_A_CTRL_PC31DOWNTO12_intermed_6 <= RIN_A_CTRL_PC31DOWNTO12_intermed_5;
		RIN_E_CTRL_PC31DOWNTO12_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 12 );
		RIN_E_CTRL_PC31DOWNTO12_intermed_2 <= RIN_E_CTRL_PC31DOWNTO12_intermed_1;
		RIN_E_CTRL_PC31DOWNTO12_intermed_3 <= RIN_E_CTRL_PC31DOWNTO12_intermed_2;
		RIN_E_CTRL_PC31DOWNTO12_intermed_4 <= RIN_E_CTRL_PC31DOWNTO12_intermed_3;
		RIN_E_CTRL_PC31DOWNTO12_intermed_5 <= RIN_E_CTRL_PC31DOWNTO12_intermed_4;
		IRIN_ADDR31DOWNTO12_intermed_1 <= IRIN.ADDR( 31 DOWNTO 12 );
		IRIN_ADDR31DOWNTO12_intermed_2 <= IRIN_ADDR31DOWNTO12_intermed_1;
		V_X_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO12_shadow;
		V_X_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_X_CTRL_PC31DOWNTO12_shadow_intermed_2;
		EX_ADD_RES32DOWNTO332DOWNTO13_shadow_intermed_1 <= EX_ADD_RES32DOWNTO332DOWNTO13_shadow;
		XC_TRAP_ADDRESS31DOWNTO12_shadow_intermed_1 <= XC_TRAP_ADDRESS31DOWNTO12_shadow;
		RIN_M_CTRL_PC31DOWNTO12_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 12 );
		RIN_M_CTRL_PC31DOWNTO12_intermed_2 <= RIN_M_CTRL_PC31DOWNTO12_intermed_1;
		RIN_M_CTRL_PC31DOWNTO12_intermed_3 <= RIN_M_CTRL_PC31DOWNTO12_intermed_2;
		RIN_M_CTRL_PC31DOWNTO12_intermed_4 <= RIN_M_CTRL_PC31DOWNTO12_intermed_3;
		IR_ADDR31DOWNTO12_intermed_1 <= IR.ADDR( 31 DOWNTO 12 );
		R_X_CTRL_PC31DOWNTO12_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 12 );
		R_X_CTRL_PC31DOWNTO12_intermed_2 <= R_X_CTRL_PC31DOWNTO12_intermed_1;
		R_D_PC31DOWNTO12_intermed_1 <= R.D.PC( 31 DOWNTO 12 );
		R_D_PC31DOWNTO12_intermed_2 <= R_D_PC31DOWNTO12_intermed_1;
		R_D_PC31DOWNTO12_intermed_3 <= R_D_PC31DOWNTO12_intermed_2;
		R_D_PC31DOWNTO12_intermed_4 <= R_D_PC31DOWNTO12_intermed_3;
		R_D_PC31DOWNTO12_intermed_5 <= R_D_PC31DOWNTO12_intermed_4;
		R_D_PC31DOWNTO12_intermed_6 <= R_D_PC31DOWNTO12_intermed_5;
		RIN_X_CTRL_PC31DOWNTO12_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 12 );
		RIN_X_CTRL_PC31DOWNTO12_intermed_2 <= RIN_X_CTRL_PC31DOWNTO12_intermed_1;
		RIN_X_CTRL_PC31DOWNTO12_intermed_3 <= RIN_X_CTRL_PC31DOWNTO12_intermed_2;
		RIN_D_PC31DOWNTO12_intermed_1 <= RIN.D.PC( 31 DOWNTO 12 );
		RIN_D_PC31DOWNTO12_intermed_2 <= RIN_D_PC31DOWNTO12_intermed_1;
		RIN_D_PC31DOWNTO12_intermed_3 <= RIN_D_PC31DOWNTO12_intermed_2;
		RIN_D_PC31DOWNTO12_intermed_4 <= RIN_D_PC31DOWNTO12_intermed_3;
		RIN_D_PC31DOWNTO12_intermed_5 <= RIN_D_PC31DOWNTO12_intermed_4;
		RIN_D_PC31DOWNTO12_intermed_6 <= RIN_D_PC31DOWNTO12_intermed_5;
		RIN_D_PC31DOWNTO12_intermed_7 <= RIN_D_PC31DOWNTO12_intermed_6;
		VIR_ADDR31DOWNTO12_shadow_intermed_1 <= VIR_ADDR31DOWNTO12_shadow;
		VIR_ADDR31DOWNTO12_shadow_intermed_2 <= VIR_ADDR31DOWNTO12_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO12_shadow;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_4 <= V_M_CTRL_PC31DOWNTO12_shadow_intermed_3;
		V_X_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_X_CTRL_TT3DOWNTO0_shadow;
		R_M_CTRL_TT3DOWNTO0_intermed_1 <= R.M.CTRL.TT( 3 DOWNTO 0 );
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1;
		R_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= R.X.RESULT( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		R_A_CTRL_TT3DOWNTO0_intermed_1 <= R.A.CTRL.TT( 3 DOWNTO 0 );
		R_A_CTRL_TT3DOWNTO0_intermed_2 <= R_A_CTRL_TT3DOWNTO0_intermed_1;
		R_A_CTRL_TT3DOWNTO0_intermed_3 <= R_A_CTRL_TT3DOWNTO0_intermed_2;
		RIN_A_CTRL_TT3DOWNTO0_intermed_1 <= RIN.A.CTRL.TT( 3 DOWNTO 0 );
		RIN_A_CTRL_TT3DOWNTO0_intermed_2 <= RIN_A_CTRL_TT3DOWNTO0_intermed_1;
		RIN_A_CTRL_TT3DOWNTO0_intermed_3 <= RIN_A_CTRL_TT3DOWNTO0_intermed_2;
		RIN_A_CTRL_TT3DOWNTO0_intermed_4 <= RIN_A_CTRL_TT3DOWNTO0_intermed_3;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_A_CTRL_TT3DOWNTO0_shadow;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_1;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_3 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_2;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_4 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_3;
		R_E_CTRL_TT3DOWNTO0_intermed_1 <= R.E.CTRL.TT( 3 DOWNTO 0 );
		R_E_CTRL_TT3DOWNTO0_intermed_2 <= R_E_CTRL_TT3DOWNTO0_intermed_1;
		RIN_M_CTRL_TT3DOWNTO0_intermed_1 <= RIN.M.CTRL.TT( 3 DOWNTO 0 );
		RIN_M_CTRL_TT3DOWNTO0_intermed_2 <= RIN_M_CTRL_TT3DOWNTO0_intermed_1;
		V_M_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_M_CTRL_TT3DOWNTO0_shadow;
		V_M_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_M_CTRL_TT3DOWNTO0_shadow_intermed_1;
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= RIN.X.RESULT( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2 <= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1;
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= RIN.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_E_CTRL_TT3DOWNTO0_shadow;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_E_CTRL_TT3DOWNTO0_shadow_intermed_1;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_3 <= V_E_CTRL_TT3DOWNTO0_shadow_intermed_2;
		RIN_X_CTRL_TT3DOWNTO0_intermed_1 <= RIN.X.CTRL.TT( 3 DOWNTO 0 );
		RIN_E_CTRL_TT3DOWNTO0_intermed_1 <= RIN.E.CTRL.TT( 3 DOWNTO 0 );
		RIN_E_CTRL_TT3DOWNTO0_intermed_2 <= RIN_E_CTRL_TT3DOWNTO0_intermed_1;
		RIN_E_CTRL_TT3DOWNTO0_intermed_3 <= RIN_E_CTRL_TT3DOWNTO0_intermed_2;
		V_X_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_X_CTRL_TT3DOWNTO0_shadow;
		V_X_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_X_CTRL_TT3DOWNTO0_shadow_intermed_1;
		R_M_CTRL_TT3DOWNTO0_intermed_1 <= R.M.CTRL.TT( 3 DOWNTO 0 );
		R_M_CTRL_TT3DOWNTO0_intermed_2 <= R_M_CTRL_TT3DOWNTO0_intermed_1;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_3 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2;
		R_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= R.X.RESULT( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		R_X_RESULT6DOWNTO03DOWNTO0_intermed_2 <= R_X_RESULT6DOWNTO03DOWNTO0_intermed_1;
		R_A_CTRL_TT3DOWNTO0_intermed_1 <= R.A.CTRL.TT( 3 DOWNTO 0 );
		R_A_CTRL_TT3DOWNTO0_intermed_2 <= R_A_CTRL_TT3DOWNTO0_intermed_1;
		R_A_CTRL_TT3DOWNTO0_intermed_3 <= R_A_CTRL_TT3DOWNTO0_intermed_2;
		R_A_CTRL_TT3DOWNTO0_intermed_4 <= R_A_CTRL_TT3DOWNTO0_intermed_3;
		RIN_A_CTRL_TT3DOWNTO0_intermed_1 <= RIN.A.CTRL.TT( 3 DOWNTO 0 );
		RIN_A_CTRL_TT3DOWNTO0_intermed_2 <= RIN_A_CTRL_TT3DOWNTO0_intermed_1;
		RIN_A_CTRL_TT3DOWNTO0_intermed_3 <= RIN_A_CTRL_TT3DOWNTO0_intermed_2;
		RIN_A_CTRL_TT3DOWNTO0_intermed_4 <= RIN_A_CTRL_TT3DOWNTO0_intermed_3;
		RIN_A_CTRL_TT3DOWNTO0_intermed_5 <= RIN_A_CTRL_TT3DOWNTO0_intermed_4;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_A_CTRL_TT3DOWNTO0_shadow;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_1;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_3 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_2;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_4 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_3;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_5 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_4;
		R_E_CTRL_TT3DOWNTO0_intermed_1 <= R.E.CTRL.TT( 3 DOWNTO 0 );
		R_E_CTRL_TT3DOWNTO0_intermed_2 <= R_E_CTRL_TT3DOWNTO0_intermed_1;
		R_E_CTRL_TT3DOWNTO0_intermed_3 <= R_E_CTRL_TT3DOWNTO0_intermed_2;
		RIN_W_S_TT3DOWNTO0_intermed_1 <= RIN.W.S.TT( 3 DOWNTO 0 );
		RIN_M_CTRL_TT3DOWNTO0_intermed_1 <= RIN.M.CTRL.TT( 3 DOWNTO 0 );
		RIN_M_CTRL_TT3DOWNTO0_intermed_2 <= RIN_M_CTRL_TT3DOWNTO0_intermed_1;
		RIN_M_CTRL_TT3DOWNTO0_intermed_3 <= RIN_M_CTRL_TT3DOWNTO0_intermed_2;
		V_M_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_M_CTRL_TT3DOWNTO0_shadow;
		V_M_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_M_CTRL_TT3DOWNTO0_shadow_intermed_1;
		V_M_CTRL_TT3DOWNTO0_shadow_intermed_3 <= V_M_CTRL_TT3DOWNTO0_shadow_intermed_2;
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= RIN.X.RESULT( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2 <= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1;
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_3 <= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2;
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= RIN.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2 <= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1;
		R_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= R.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_E_CTRL_TT3DOWNTO0_shadow;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_E_CTRL_TT3DOWNTO0_shadow_intermed_1;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_3 <= V_E_CTRL_TT3DOWNTO0_shadow_intermed_2;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_4 <= V_E_CTRL_TT3DOWNTO0_shadow_intermed_3;
		RIN_X_CTRL_TT3DOWNTO0_intermed_1 <= RIN.X.CTRL.TT( 3 DOWNTO 0 );
		RIN_X_CTRL_TT3DOWNTO0_intermed_2 <= RIN_X_CTRL_TT3DOWNTO0_intermed_1;
		R_X_CTRL_TT3DOWNTO0_intermed_1 <= R.X.CTRL.TT( 3 DOWNTO 0 );
		RIN_E_CTRL_TT3DOWNTO0_intermed_1 <= RIN.E.CTRL.TT( 3 DOWNTO 0 );
		RIN_E_CTRL_TT3DOWNTO0_intermed_2 <= RIN_E_CTRL_TT3DOWNTO0_intermed_1;
		RIN_E_CTRL_TT3DOWNTO0_intermed_3 <= RIN_E_CTRL_TT3DOWNTO0_intermed_2;
		RIN_E_CTRL_TT3DOWNTO0_intermed_4 <= RIN_E_CTRL_TT3DOWNTO0_intermed_3;
		XC_VECTT3DOWNTO0_shadow_intermed_1 <= XC_VECTT3DOWNTO0_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		V_X_DATA03_shadow_intermed_1 <= V_X_DATA03_shadow;
		V_X_DATA03_shadow_intermed_2 <= V_X_DATA03_shadow_intermed_1;
		DCO_DATA03_intermed_1 <= DCO.DATA ( 0 )( 3 );
		RIN_X_DATA03_intermed_1 <= RIN.X.DATA ( 0 )( 3 );
		R_X_DATA03_intermed_1 <= R.X.DATA( 0 )( 3 );
		RIN_X_DATA03_intermed_1 <= RIN.X.DATA( 0 )( 3 );
		RIN_X_DATA03_intermed_2 <= RIN_X_DATA03_intermed_1;
		R_M_CTRL_PC31DOWNTO12_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 12 );
		R_M_CTRL_PC31DOWNTO12_intermed_2 <= R_M_CTRL_PC31DOWNTO12_intermed_1;
		V_D_PC31DOWNTO12_shadow_intermed_1 <= V_D_PC31DOWNTO12_shadow;
		V_D_PC31DOWNTO12_shadow_intermed_2 <= V_D_PC31DOWNTO12_shadow_intermed_1;
		V_D_PC31DOWNTO12_shadow_intermed_3 <= V_D_PC31DOWNTO12_shadow_intermed_2;
		V_D_PC31DOWNTO12_shadow_intermed_4 <= V_D_PC31DOWNTO12_shadow_intermed_3;
		V_D_PC31DOWNTO12_shadow_intermed_5 <= V_D_PC31DOWNTO12_shadow_intermed_4;
		V_D_PC31DOWNTO12_shadow_intermed_6 <= V_D_PC31DOWNTO12_shadow_intermed_5;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO12_shadow;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_4;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO12_shadow;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_3;
		R_A_CTRL_PC31DOWNTO12_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 12 );
		R_A_CTRL_PC31DOWNTO12_intermed_2 <= R_A_CTRL_PC31DOWNTO12_intermed_1;
		R_A_CTRL_PC31DOWNTO12_intermed_3 <= R_A_CTRL_PC31DOWNTO12_intermed_2;
		R_A_CTRL_PC31DOWNTO12_intermed_4 <= R_A_CTRL_PC31DOWNTO12_intermed_3;
		R_E_CTRL_PC31DOWNTO12_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 12 );
		R_E_CTRL_PC31DOWNTO12_intermed_2 <= R_E_CTRL_PC31DOWNTO12_intermed_1;
		R_E_CTRL_PC31DOWNTO12_intermed_3 <= R_E_CTRL_PC31DOWNTO12_intermed_2;
		RIN_A_CTRL_PC31DOWNTO12_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 12 );
		RIN_A_CTRL_PC31DOWNTO12_intermed_2 <= RIN_A_CTRL_PC31DOWNTO12_intermed_1;
		RIN_A_CTRL_PC31DOWNTO12_intermed_3 <= RIN_A_CTRL_PC31DOWNTO12_intermed_2;
		RIN_A_CTRL_PC31DOWNTO12_intermed_4 <= RIN_A_CTRL_PC31DOWNTO12_intermed_3;
		RIN_A_CTRL_PC31DOWNTO12_intermed_5 <= RIN_A_CTRL_PC31DOWNTO12_intermed_4;
		RIN_E_CTRL_PC31DOWNTO12_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 12 );
		RIN_E_CTRL_PC31DOWNTO12_intermed_2 <= RIN_E_CTRL_PC31DOWNTO12_intermed_1;
		RIN_E_CTRL_PC31DOWNTO12_intermed_3 <= RIN_E_CTRL_PC31DOWNTO12_intermed_2;
		RIN_E_CTRL_PC31DOWNTO12_intermed_4 <= RIN_E_CTRL_PC31DOWNTO12_intermed_3;
		IRIN_ADDR31DOWNTO12_intermed_1 <= IRIN.ADDR( 31 DOWNTO 12 );
		V_X_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO12_shadow;
		V_X_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO12_shadow_intermed_1;
		RIN_M_CTRL_PC31DOWNTO12_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 12 );
		RIN_M_CTRL_PC31DOWNTO12_intermed_2 <= RIN_M_CTRL_PC31DOWNTO12_intermed_1;
		RIN_M_CTRL_PC31DOWNTO12_intermed_3 <= RIN_M_CTRL_PC31DOWNTO12_intermed_2;
		R_X_CTRL_PC31DOWNTO12_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 12 );
		R_D_PC31DOWNTO12_intermed_1 <= R.D.PC( 31 DOWNTO 12 );
		R_D_PC31DOWNTO12_intermed_2 <= R_D_PC31DOWNTO12_intermed_1;
		R_D_PC31DOWNTO12_intermed_3 <= R_D_PC31DOWNTO12_intermed_2;
		R_D_PC31DOWNTO12_intermed_4 <= R_D_PC31DOWNTO12_intermed_3;
		R_D_PC31DOWNTO12_intermed_5 <= R_D_PC31DOWNTO12_intermed_4;
		RIN_X_CTRL_PC31DOWNTO12_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 12 );
		RIN_X_CTRL_PC31DOWNTO12_intermed_2 <= RIN_X_CTRL_PC31DOWNTO12_intermed_1;
		RIN_D_PC31DOWNTO12_intermed_1 <= RIN.D.PC( 31 DOWNTO 12 );
		RIN_D_PC31DOWNTO12_intermed_2 <= RIN_D_PC31DOWNTO12_intermed_1;
		RIN_D_PC31DOWNTO12_intermed_3 <= RIN_D_PC31DOWNTO12_intermed_2;
		RIN_D_PC31DOWNTO12_intermed_4 <= RIN_D_PC31DOWNTO12_intermed_3;
		RIN_D_PC31DOWNTO12_intermed_5 <= RIN_D_PC31DOWNTO12_intermed_4;
		RIN_D_PC31DOWNTO12_intermed_6 <= RIN_D_PC31DOWNTO12_intermed_5;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO12_shadow;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO12_shadow_intermed_2;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		RIN_M_CTRL_PC31DOWNTO2_intermed_2 <= RIN_M_CTRL_PC31DOWNTO2_intermed_1;
		RIN_M_CTRL_PC31DOWNTO2_intermed_3 <= RIN_M_CTRL_PC31DOWNTO2_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		V_D_PC31DOWNTO2_shadow_intermed_5 <= V_D_PC31DOWNTO2_shadow_intermed_4;
		V_D_PC31DOWNTO2_shadow_intermed_6 <= V_D_PC31DOWNTO2_shadow_intermed_5;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_5 <= RIN_D_PC31DOWNTO2_intermed_4;
		RIN_D_PC31DOWNTO2_intermed_6 <= RIN_D_PC31DOWNTO2_intermed_5;
		RIN_X_CTRL_PC31DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 2 );
		RIN_X_CTRL_PC31DOWNTO2_intermed_2 <= RIN_X_CTRL_PC31DOWNTO2_intermed_1;
		IRIN_ADDR31DOWNTO2_intermed_1 <= IRIN.ADDR( 31 DOWNTO 2 );
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		R_D_PC31DOWNTO2_intermed_4 <= R_D_PC31DOWNTO2_intermed_3;
		R_D_PC31DOWNTO2_intermed_5 <= R_D_PC31DOWNTO2_intermed_4;
		R_M_CTRL_PC31DOWNTO2_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 2 );
		R_M_CTRL_PC31DOWNTO2_intermed_2 <= R_M_CTRL_PC31DOWNTO2_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		RIN_A_CTRL_PC31DOWNTO2_intermed_4 <= RIN_A_CTRL_PC31DOWNTO2_intermed_3;
		RIN_A_CTRL_PC31DOWNTO2_intermed_5 <= RIN_A_CTRL_PC31DOWNTO2_intermed_4;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_3 <= R_A_CTRL_PC31DOWNTO2_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_4 <= R_A_CTRL_PC31DOWNTO2_intermed_3;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO2_shadow;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2;
		R_X_CTRL_PC31DOWNTO2_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		R_E_CTRL_PC31DOWNTO2_intermed_2 <= R_E_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_3 <= R_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_E_CTRL_PC31DOWNTO2_intermed_3 <= RIN_E_CTRL_PC31DOWNTO2_intermed_2;
		RIN_E_CTRL_PC31DOWNTO2_intermed_4 <= RIN_E_CTRL_PC31DOWNTO2_intermed_3;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO2_shadow;
		V_X_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_F_PC31DOWNTO4_shadow_intermed_1 <= V_F_PC31DOWNTO4_shadow;
		V_X_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_X_CTRL_PC31DOWNTO4_shadow;
		V_X_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_X_CTRL_PC31DOWNTO4_shadow_intermed_1;
		V_X_CTRL_PC31DOWNTO4_shadow_intermed_3 <= V_X_CTRL_PC31DOWNTO4_shadow_intermed_2;
		IR_ADDR31DOWNTO4_intermed_1 <= IR.ADDR( 31 DOWNTO 4 );
		VIR_ADDR31DOWNTO4_shadow_intermed_1 <= VIR_ADDR31DOWNTO4_shadow;
		VIR_ADDR31DOWNTO4_shadow_intermed_2 <= VIR_ADDR31DOWNTO4_shadow_intermed_1;
		RIN_F_PC31DOWNTO4_intermed_1 <= RIN.F.PC( 31 DOWNTO 4 );
		RIN_A_CTRL_PC31DOWNTO4_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 4 );
		RIN_A_CTRL_PC31DOWNTO4_intermed_2 <= RIN_A_CTRL_PC31DOWNTO4_intermed_1;
		RIN_A_CTRL_PC31DOWNTO4_intermed_3 <= RIN_A_CTRL_PC31DOWNTO4_intermed_2;
		RIN_A_CTRL_PC31DOWNTO4_intermed_4 <= RIN_A_CTRL_PC31DOWNTO4_intermed_3;
		RIN_A_CTRL_PC31DOWNTO4_intermed_5 <= RIN_A_CTRL_PC31DOWNTO4_intermed_4;
		RIN_A_CTRL_PC31DOWNTO4_intermed_6 <= RIN_A_CTRL_PC31DOWNTO4_intermed_5;
		R_A_CTRL_PC31DOWNTO4_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 4 );
		R_A_CTRL_PC31DOWNTO4_intermed_2 <= R_A_CTRL_PC31DOWNTO4_intermed_1;
		R_A_CTRL_PC31DOWNTO4_intermed_3 <= R_A_CTRL_PC31DOWNTO4_intermed_2;
		R_A_CTRL_PC31DOWNTO4_intermed_4 <= R_A_CTRL_PC31DOWNTO4_intermed_3;
		R_A_CTRL_PC31DOWNTO4_intermed_5 <= R_A_CTRL_PC31DOWNTO4_intermed_4;
		R_D_PC31DOWNTO4_intermed_1 <= R.D.PC( 31 DOWNTO 4 );
		R_D_PC31DOWNTO4_intermed_2 <= R_D_PC31DOWNTO4_intermed_1;
		R_D_PC31DOWNTO4_intermed_3 <= R_D_PC31DOWNTO4_intermed_2;
		R_D_PC31DOWNTO4_intermed_4 <= R_D_PC31DOWNTO4_intermed_3;
		R_D_PC31DOWNTO4_intermed_5 <= R_D_PC31DOWNTO4_intermed_4;
		R_D_PC31DOWNTO4_intermed_6 <= R_D_PC31DOWNTO4_intermed_5;
		RIN_X_CTRL_PC31DOWNTO4_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 4 );
		RIN_X_CTRL_PC31DOWNTO4_intermed_2 <= RIN_X_CTRL_PC31DOWNTO4_intermed_1;
		RIN_X_CTRL_PC31DOWNTO4_intermed_3 <= RIN_X_CTRL_PC31DOWNTO4_intermed_2;
		EX_ADD_RES32DOWNTO332DOWNTO5_shadow_intermed_1 <= EX_ADD_RES32DOWNTO332DOWNTO5_shadow;
		V_D_PC31DOWNTO4_shadow_intermed_1 <= V_D_PC31DOWNTO4_shadow;
		V_D_PC31DOWNTO4_shadow_intermed_2 <= V_D_PC31DOWNTO4_shadow_intermed_1;
		V_D_PC31DOWNTO4_shadow_intermed_3 <= V_D_PC31DOWNTO4_shadow_intermed_2;
		V_D_PC31DOWNTO4_shadow_intermed_4 <= V_D_PC31DOWNTO4_shadow_intermed_3;
		V_D_PC31DOWNTO4_shadow_intermed_5 <= V_D_PC31DOWNTO4_shadow_intermed_4;
		V_D_PC31DOWNTO4_shadow_intermed_6 <= V_D_PC31DOWNTO4_shadow_intermed_5;
		V_D_PC31DOWNTO4_shadow_intermed_7 <= V_D_PC31DOWNTO4_shadow_intermed_6;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO4_shadow;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO4_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO4_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_4 <= V_E_CTRL_PC31DOWNTO4_shadow_intermed_3;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_5 <= V_E_CTRL_PC31DOWNTO4_shadow_intermed_4;
		RIN_M_CTRL_PC31DOWNTO4_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 4 );
		RIN_M_CTRL_PC31DOWNTO4_intermed_2 <= RIN_M_CTRL_PC31DOWNTO4_intermed_1;
		RIN_M_CTRL_PC31DOWNTO4_intermed_3 <= RIN_M_CTRL_PC31DOWNTO4_intermed_2;
		RIN_M_CTRL_PC31DOWNTO4_intermed_4 <= RIN_M_CTRL_PC31DOWNTO4_intermed_3;
		R_X_CTRL_PC31DOWNTO4_intermed_1 <= R.X.CTRL.PC( 31 DOWNTO 4 );
		R_X_CTRL_PC31DOWNTO4_intermed_2 <= R_X_CTRL_PC31DOWNTO4_intermed_1;
		IRIN_ADDR31DOWNTO4_intermed_1 <= IRIN.ADDR( 31 DOWNTO 4 );
		IRIN_ADDR31DOWNTO4_intermed_2 <= IRIN_ADDR31DOWNTO4_intermed_1;
		V_M_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO4_shadow;
		V_M_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO4_shadow_intermed_1;
		V_M_CTRL_PC31DOWNTO4_shadow_intermed_3 <= V_M_CTRL_PC31DOWNTO4_shadow_intermed_2;
		V_M_CTRL_PC31DOWNTO4_shadow_intermed_4 <= V_M_CTRL_PC31DOWNTO4_shadow_intermed_3;
		R_M_CTRL_PC31DOWNTO4_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 4 );
		R_M_CTRL_PC31DOWNTO4_intermed_2 <= R_M_CTRL_PC31DOWNTO4_intermed_1;
		R_M_CTRL_PC31DOWNTO4_intermed_3 <= R_M_CTRL_PC31DOWNTO4_intermed_2;
		RIN_D_PC31DOWNTO4_intermed_1 <= RIN.D.PC( 31 DOWNTO 4 );
		RIN_D_PC31DOWNTO4_intermed_2 <= RIN_D_PC31DOWNTO4_intermed_1;
		RIN_D_PC31DOWNTO4_intermed_3 <= RIN_D_PC31DOWNTO4_intermed_2;
		RIN_D_PC31DOWNTO4_intermed_4 <= RIN_D_PC31DOWNTO4_intermed_3;
		RIN_D_PC31DOWNTO4_intermed_5 <= RIN_D_PC31DOWNTO4_intermed_4;
		RIN_D_PC31DOWNTO4_intermed_6 <= RIN_D_PC31DOWNTO4_intermed_5;
		RIN_D_PC31DOWNTO4_intermed_7 <= RIN_D_PC31DOWNTO4_intermed_6;
		RIN_E_CTRL_PC31DOWNTO4_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 4 );
		RIN_E_CTRL_PC31DOWNTO4_intermed_2 <= RIN_E_CTRL_PC31DOWNTO4_intermed_1;
		RIN_E_CTRL_PC31DOWNTO4_intermed_3 <= RIN_E_CTRL_PC31DOWNTO4_intermed_2;
		RIN_E_CTRL_PC31DOWNTO4_intermed_4 <= RIN_E_CTRL_PC31DOWNTO4_intermed_3;
		RIN_E_CTRL_PC31DOWNTO4_intermed_5 <= RIN_E_CTRL_PC31DOWNTO4_intermed_4;
		EX_JUMP_ADDRESS31DOWNTO4_shadow_intermed_1 <= EX_JUMP_ADDRESS31DOWNTO4_shadow;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO4_shadow;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_5 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_4;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_6 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_5;
		R_E_CTRL_PC31DOWNTO4_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 4 );
		R_E_CTRL_PC31DOWNTO4_intermed_2 <= R_E_CTRL_PC31DOWNTO4_intermed_1;
		R_E_CTRL_PC31DOWNTO4_intermed_3 <= R_E_CTRL_PC31DOWNTO4_intermed_2;
		R_E_CTRL_PC31DOWNTO4_intermed_4 <= R_E_CTRL_PC31DOWNTO4_intermed_3;
		R_D_PC3DOWNTO2_intermed_1 <= R.D.PC( 3 DOWNTO 2 );
		R_D_PC3DOWNTO2_intermed_2 <= R_D_PC3DOWNTO2_intermed_1;
		R_D_PC3DOWNTO2_intermed_3 <= R_D_PC3DOWNTO2_intermed_2;
		R_D_PC3DOWNTO2_intermed_4 <= R_D_PC3DOWNTO2_intermed_3;
		R_D_PC3DOWNTO2_intermed_5 <= R_D_PC3DOWNTO2_intermed_4;
		R_D_PC3DOWNTO2_intermed_6 <= R_D_PC3DOWNTO2_intermed_5;
		V_D_PC3DOWNTO2_shadow_intermed_1 <= V_D_PC3DOWNTO2_shadow;
		V_D_PC3DOWNTO2_shadow_intermed_2 <= V_D_PC3DOWNTO2_shadow_intermed_1;
		V_D_PC3DOWNTO2_shadow_intermed_3 <= V_D_PC3DOWNTO2_shadow_intermed_2;
		V_D_PC3DOWNTO2_shadow_intermed_4 <= V_D_PC3DOWNTO2_shadow_intermed_3;
		V_D_PC3DOWNTO2_shadow_intermed_5 <= V_D_PC3DOWNTO2_shadow_intermed_4;
		V_D_PC3DOWNTO2_shadow_intermed_6 <= V_D_PC3DOWNTO2_shadow_intermed_5;
		V_D_PC3DOWNTO2_shadow_intermed_7 <= V_D_PC3DOWNTO2_shadow_intermed_6;
		VIR_ADDR3DOWNTO2_shadow_intermed_1 <= VIR_ADDR3DOWNTO2_shadow;
		VIR_ADDR3DOWNTO2_shadow_intermed_2 <= VIR_ADDR3DOWNTO2_shadow_intermed_1;
		RIN_D_PC3DOWNTO2_intermed_1 <= RIN.D.PC( 3 DOWNTO 2 );
		RIN_D_PC3DOWNTO2_intermed_2 <= RIN_D_PC3DOWNTO2_intermed_1;
		RIN_D_PC3DOWNTO2_intermed_3 <= RIN_D_PC3DOWNTO2_intermed_2;
		RIN_D_PC3DOWNTO2_intermed_4 <= RIN_D_PC3DOWNTO2_intermed_3;
		RIN_D_PC3DOWNTO2_intermed_5 <= RIN_D_PC3DOWNTO2_intermed_4;
		RIN_D_PC3DOWNTO2_intermed_6 <= RIN_D_PC3DOWNTO2_intermed_5;
		RIN_D_PC3DOWNTO2_intermed_7 <= RIN_D_PC3DOWNTO2_intermed_6;
		R_M_CTRL_PC3DOWNTO2_intermed_1 <= R.M.CTRL.PC( 3 DOWNTO 2 );
		R_M_CTRL_PC3DOWNTO2_intermed_2 <= R_M_CTRL_PC3DOWNTO2_intermed_1;
		R_M_CTRL_PC3DOWNTO2_intermed_3 <= R_M_CTRL_PC3DOWNTO2_intermed_2;
		R_E_CTRL_PC3DOWNTO2_intermed_1 <= R.E.CTRL.PC( 3 DOWNTO 2 );
		R_E_CTRL_PC3DOWNTO2_intermed_2 <= R_E_CTRL_PC3DOWNTO2_intermed_1;
		R_E_CTRL_PC3DOWNTO2_intermed_3 <= R_E_CTRL_PC3DOWNTO2_intermed_2;
		R_E_CTRL_PC3DOWNTO2_intermed_4 <= R_E_CTRL_PC3DOWNTO2_intermed_3;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC3DOWNTO2_shadow;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC3DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC3DOWNTO2_shadow_intermed_2;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_4 <= V_E_CTRL_PC3DOWNTO2_shadow_intermed_3;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_5 <= V_E_CTRL_PC3DOWNTO2_shadow_intermed_4;
		RIN_X_CTRL_PC3DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 3 DOWNTO 2 );
		RIN_X_CTRL_PC3DOWNTO2_intermed_2 <= RIN_X_CTRL_PC3DOWNTO2_intermed_1;
		RIN_X_CTRL_PC3DOWNTO2_intermed_3 <= RIN_X_CTRL_PC3DOWNTO2_intermed_2;
		R_A_CTRL_PC3DOWNTO2_intermed_1 <= R.A.CTRL.PC( 3 DOWNTO 2 );
		R_A_CTRL_PC3DOWNTO2_intermed_2 <= R_A_CTRL_PC3DOWNTO2_intermed_1;
		R_A_CTRL_PC3DOWNTO2_intermed_3 <= R_A_CTRL_PC3DOWNTO2_intermed_2;
		R_A_CTRL_PC3DOWNTO2_intermed_4 <= R_A_CTRL_PC3DOWNTO2_intermed_3;
		R_A_CTRL_PC3DOWNTO2_intermed_5 <= R_A_CTRL_PC3DOWNTO2_intermed_4;
		V_X_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_X_CTRL_PC3DOWNTO2_shadow;
		V_X_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_X_CTRL_PC3DOWNTO2_shadow_intermed_1;
		V_X_CTRL_PC3DOWNTO2_shadow_intermed_3 <= V_X_CTRL_PC3DOWNTO2_shadow_intermed_2;
		RIN_M_CTRL_PC3DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 3 DOWNTO 2 );
		RIN_M_CTRL_PC3DOWNTO2_intermed_2 <= RIN_M_CTRL_PC3DOWNTO2_intermed_1;
		RIN_M_CTRL_PC3DOWNTO2_intermed_3 <= RIN_M_CTRL_PC3DOWNTO2_intermed_2;
		RIN_M_CTRL_PC3DOWNTO2_intermed_4 <= RIN_M_CTRL_PC3DOWNTO2_intermed_3;
		IRIN_ADDR3DOWNTO2_intermed_1 <= IRIN.ADDR( 3 DOWNTO 2 );
		IRIN_ADDR3DOWNTO2_intermed_2 <= IRIN_ADDR3DOWNTO2_intermed_1;
		EX_JUMP_ADDRESS3DOWNTO2_shadow_intermed_1 <= EX_JUMP_ADDRESS3DOWNTO2_shadow;
		EX_ADD_RES32DOWNTO34DOWNTO3_shadow_intermed_1 <= EX_ADD_RES32DOWNTO34DOWNTO3_shadow;
		RIN_A_CTRL_PC3DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 3 DOWNTO 2 );
		RIN_A_CTRL_PC3DOWNTO2_intermed_2 <= RIN_A_CTRL_PC3DOWNTO2_intermed_1;
		RIN_A_CTRL_PC3DOWNTO2_intermed_3 <= RIN_A_CTRL_PC3DOWNTO2_intermed_2;
		RIN_A_CTRL_PC3DOWNTO2_intermed_4 <= RIN_A_CTRL_PC3DOWNTO2_intermed_3;
		RIN_A_CTRL_PC3DOWNTO2_intermed_5 <= RIN_A_CTRL_PC3DOWNTO2_intermed_4;
		RIN_A_CTRL_PC3DOWNTO2_intermed_6 <= RIN_A_CTRL_PC3DOWNTO2_intermed_5;
		V_F_PC3DOWNTO2_shadow_intermed_1 <= V_F_PC3DOWNTO2_shadow;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC3DOWNTO2_shadow;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_3;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_5 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_4;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_6 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_5;
		IR_ADDR3DOWNTO2_intermed_1 <= IR.ADDR( 3 DOWNTO 2 );
		V_M_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC3DOWNTO2_shadow;
		V_M_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC3DOWNTO2_shadow_intermed_1;
		V_M_CTRL_PC3DOWNTO2_shadow_intermed_3 <= V_M_CTRL_PC3DOWNTO2_shadow_intermed_2;
		V_M_CTRL_PC3DOWNTO2_shadow_intermed_4 <= V_M_CTRL_PC3DOWNTO2_shadow_intermed_3;
		R_X_CTRL_PC3DOWNTO2_intermed_1 <= R.X.CTRL.PC( 3 DOWNTO 2 );
		R_X_CTRL_PC3DOWNTO2_intermed_2 <= R_X_CTRL_PC3DOWNTO2_intermed_1;
		RIN_E_CTRL_PC3DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 3 DOWNTO 2 );
		RIN_E_CTRL_PC3DOWNTO2_intermed_2 <= RIN_E_CTRL_PC3DOWNTO2_intermed_1;
		RIN_E_CTRL_PC3DOWNTO2_intermed_3 <= RIN_E_CTRL_PC3DOWNTO2_intermed_2;
		RIN_E_CTRL_PC3DOWNTO2_intermed_4 <= RIN_E_CTRL_PC3DOWNTO2_intermed_3;
		RIN_E_CTRL_PC3DOWNTO2_intermed_5 <= RIN_E_CTRL_PC3DOWNTO2_intermed_4;
		RIN_F_PC3DOWNTO2_intermed_1 <= RIN.F.PC( 3 DOWNTO 2 );
		V_E_CTRL_RD7DOWNTO0_shadow_intermed_1 <= V_E_CTRL_RD7DOWNTO0_shadow;
		V_E_CTRL_RD7DOWNTO0_shadow_intermed_2 <= V_E_CTRL_RD7DOWNTO0_shadow_intermed_1;
		R_E_CTRL_RD7DOWNTO0_intermed_1 <= R.E.CTRL.RD ( 7 DOWNTO 0 );
		V_A_CTRL_RD7DOWNTO0_shadow_intermed_1 <= V_A_CTRL_RD7DOWNTO0_shadow;
		V_A_CTRL_RD7DOWNTO0_shadow_intermed_2 <= V_A_CTRL_RD7DOWNTO0_shadow_intermed_1;
		V_A_CTRL_RD7DOWNTO0_shadow_intermed_3 <= V_A_CTRL_RD7DOWNTO0_shadow_intermed_2;
		RIN_A_CTRL_RD7DOWNTO0_intermed_1 <= RIN.A.CTRL.RD ( 7 DOWNTO 0 );
		RIN_A_CTRL_RD7DOWNTO0_intermed_2 <= RIN_A_CTRL_RD7DOWNTO0_intermed_1;
		RIN_A_CTRL_RD7DOWNTO0_intermed_3 <= RIN_A_CTRL_RD7DOWNTO0_intermed_2;
		R_A_CTRL_RD7DOWNTO0_intermed_1 <= R.A.CTRL.RD ( 7 DOWNTO 0 );
		R_A_CTRL_RD7DOWNTO0_intermed_2 <= R_A_CTRL_RD7DOWNTO0_intermed_1;
		RIN_E_CTRL_RD7DOWNTO0_intermed_1 <= RIN.E.CTRL.RD ( 7 DOWNTO 0 );
		RIN_E_CTRL_RD7DOWNTO0_intermed_2 <= RIN_E_CTRL_RD7DOWNTO0_intermed_1;
		RIN_M_CTRL_RD7DOWNTO0_intermed_1 <= RIN.M.CTRL.RD ( 7 DOWNTO 0 );
		RIN_D_PC_intermed_1 <= RIN.D.PC;
		RIN_D_PC_intermed_2 <= RIN_D_PC_intermed_1;
		RIN_D_PC_intermed_3 <= RIN_D_PC_intermed_2;
		RIN_D_PC_intermed_4 <= RIN_D_PC_intermed_3;
		RIN_A_CTRL_PC_intermed_1 <= RIN.A.CTRL.PC;
		RIN_A_CTRL_PC_intermed_2 <= RIN_A_CTRL_PC_intermed_1;
		RIN_A_CTRL_PC_intermed_3 <= RIN_A_CTRL_PC_intermed_2;
		R_A_CTRL_PC_intermed_1 <= R.A.CTRL.PC;
		R_A_CTRL_PC_intermed_2 <= R_A_CTRL_PC_intermed_1;
		V_E_CTRL_PC_shadow_intermed_1 <= V_E_CTRL_PC_shadow;
		V_E_CTRL_PC_shadow_intermed_2 <= V_E_CTRL_PC_shadow_intermed_1;
		R_E_CTRL_PC_intermed_1 <= R.E.CTRL.PC;
		RIN_M_CTRL_PC_intermed_1 <= RIN.M.CTRL.PC;
		V_A_CTRL_PC_shadow_intermed_1 <= V_A_CTRL_PC_shadow;
		V_A_CTRL_PC_shadow_intermed_2 <= V_A_CTRL_PC_shadow_intermed_1;
		V_A_CTRL_PC_shadow_intermed_3 <= V_A_CTRL_PC_shadow_intermed_2;
		R_D_PC_intermed_1 <= R.D.PC;
		R_D_PC_intermed_2 <= R_D_PC_intermed_1;
		R_D_PC_intermed_3 <= R_D_PC_intermed_2;
		RIN_E_CTRL_PC_intermed_1 <= RIN.E.CTRL.PC;
		RIN_E_CTRL_PC_intermed_2 <= RIN_E_CTRL_PC_intermed_1;
		V_D_PC_shadow_intermed_1 <= V_D_PC_shadow;
		V_D_PC_shadow_intermed_2 <= V_D_PC_shadow_intermed_1;
		V_D_PC_shadow_intermed_3 <= V_D_PC_shadow_intermed_2;
		V_D_PC_shadow_intermed_4 <= V_D_PC_shadow_intermed_3;
		RIN_M_CTRL_PC31DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 2 );
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_4 <= V_D_PC31DOWNTO2_shadow_intermed_3;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_4 <= RIN_D_PC31DOWNTO2_intermed_3;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		R_D_PC31DOWNTO2_intermed_3 <= R_D_PC31DOWNTO2_intermed_2;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO2_shadow;
		V_E_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_3 <= RIN_A_CTRL_PC31DOWNTO2_intermed_2;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		R_A_CTRL_PC31DOWNTO2_intermed_2 <= R_A_CTRL_PC31DOWNTO2_intermed_1;
		R_E_CTRL_PC31DOWNTO2_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_2 <= RIN_E_CTRL_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_INST20_intermed_1 <= RIN.A.CTRL.INST ( 20 );
		RIN_A_CTRL_INST20_intermed_1 <= RIN.A.CTRL.INST( 20 );
		RIN_A_CTRL_INST20_intermed_2 <= RIN_A_CTRL_INST20_intermed_1;
		V_A_CTRL_INST20_shadow_intermed_1 <= V_A_CTRL_INST20_shadow;
		V_A_CTRL_INST20_shadow_intermed_2 <= V_A_CTRL_INST20_shadow_intermed_1;
		DE_INST20_shadow_intermed_1 <= DE_INST20_shadow;
		R_A_CTRL_INST20_intermed_1 <= R.A.CTRL.INST( 20 );
		RIN_A_CTRL_INST20_intermed_1 <= RIN.A.CTRL.INST( 20 );
		DE_INST20_shadow_intermed_1 <= DE_INST20_shadow;
		R_A_CTRL_INST24_intermed_1 <= R.A.CTRL.INST( 24 );
		RIN_A_CTRL_INST24_intermed_1 <= RIN.A.CTRL.INST( 24 );
		RIN_A_CTRL_INST24_intermed_2 <= RIN_A_CTRL_INST24_intermed_1;
		V_A_CTRL_INST24_shadow_intermed_1 <= V_A_CTRL_INST24_shadow;
		V_A_CTRL_INST24_shadow_intermed_2 <= V_A_CTRL_INST24_shadow_intermed_1;
		DE_INST24_shadow_intermed_1 <= DE_INST24_shadow;
		RIN_A_CTRL_INST24_intermed_1 <= RIN.A.CTRL.INST ( 24 );
		RIN_A_CTRL_INST24_intermed_1 <= RIN.A.CTRL.INST( 24 );
		DE_INST24_shadow_intermed_1 <= DE_INST24_shadow;
		RIN_A_CTRL_PC31DOWNTO4_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 4 );
		RIN_A_CTRL_PC31DOWNTO4_intermed_2 <= RIN_A_CTRL_PC31DOWNTO4_intermed_1;
		RIN_A_CTRL_PC31DOWNTO4_intermed_3 <= RIN_A_CTRL_PC31DOWNTO4_intermed_2;
		RIN_A_CTRL_PC31DOWNTO4_intermed_4 <= RIN_A_CTRL_PC31DOWNTO4_intermed_3;
		R_A_CTRL_PC31DOWNTO4_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 4 );
		R_A_CTRL_PC31DOWNTO4_intermed_2 <= R_A_CTRL_PC31DOWNTO4_intermed_1;
		R_A_CTRL_PC31DOWNTO4_intermed_3 <= R_A_CTRL_PC31DOWNTO4_intermed_2;
		R_D_PC31DOWNTO4_intermed_1 <= R.D.PC( 31 DOWNTO 4 );
		R_D_PC31DOWNTO4_intermed_2 <= R_D_PC31DOWNTO4_intermed_1;
		R_D_PC31DOWNTO4_intermed_3 <= R_D_PC31DOWNTO4_intermed_2;
		R_D_PC31DOWNTO4_intermed_4 <= R_D_PC31DOWNTO4_intermed_3;
		RIN_X_CTRL_PC31DOWNTO4_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 4 );
		V_D_PC31DOWNTO4_shadow_intermed_1 <= V_D_PC31DOWNTO4_shadow;
		V_D_PC31DOWNTO4_shadow_intermed_2 <= V_D_PC31DOWNTO4_shadow_intermed_1;
		V_D_PC31DOWNTO4_shadow_intermed_3 <= V_D_PC31DOWNTO4_shadow_intermed_2;
		V_D_PC31DOWNTO4_shadow_intermed_4 <= V_D_PC31DOWNTO4_shadow_intermed_3;
		V_D_PC31DOWNTO4_shadow_intermed_5 <= V_D_PC31DOWNTO4_shadow_intermed_4;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO4_shadow;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO4_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO4_shadow_intermed_2;
		RIN_M_CTRL_PC31DOWNTO4_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 4 );
		RIN_M_CTRL_PC31DOWNTO4_intermed_2 <= RIN_M_CTRL_PC31DOWNTO4_intermed_1;
		V_M_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO4_shadow;
		V_M_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO4_shadow_intermed_1;
		R_M_CTRL_PC31DOWNTO4_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 4 );
		RIN_D_PC31DOWNTO4_intermed_1 <= RIN.D.PC( 31 DOWNTO 4 );
		RIN_D_PC31DOWNTO4_intermed_2 <= RIN_D_PC31DOWNTO4_intermed_1;
		RIN_D_PC31DOWNTO4_intermed_3 <= RIN_D_PC31DOWNTO4_intermed_2;
		RIN_D_PC31DOWNTO4_intermed_4 <= RIN_D_PC31DOWNTO4_intermed_3;
		RIN_D_PC31DOWNTO4_intermed_5 <= RIN_D_PC31DOWNTO4_intermed_4;
		RIN_E_CTRL_PC31DOWNTO4_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 4 );
		RIN_E_CTRL_PC31DOWNTO4_intermed_2 <= RIN_E_CTRL_PC31DOWNTO4_intermed_1;
		RIN_E_CTRL_PC31DOWNTO4_intermed_3 <= RIN_E_CTRL_PC31DOWNTO4_intermed_2;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO4_shadow;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_3;
		R_E_CTRL_PC31DOWNTO4_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 4 );
		R_E_CTRL_PC31DOWNTO4_intermed_2 <= R_E_CTRL_PC31DOWNTO4_intermed_1;
		R_D_PC3DOWNTO2_intermed_1 <= R.D.PC( 3 DOWNTO 2 );
		R_D_PC3DOWNTO2_intermed_2 <= R_D_PC3DOWNTO2_intermed_1;
		R_D_PC3DOWNTO2_intermed_3 <= R_D_PC3DOWNTO2_intermed_2;
		R_D_PC3DOWNTO2_intermed_4 <= R_D_PC3DOWNTO2_intermed_3;
		V_D_PC3DOWNTO2_shadow_intermed_1 <= V_D_PC3DOWNTO2_shadow;
		V_D_PC3DOWNTO2_shadow_intermed_2 <= V_D_PC3DOWNTO2_shadow_intermed_1;
		V_D_PC3DOWNTO2_shadow_intermed_3 <= V_D_PC3DOWNTO2_shadow_intermed_2;
		V_D_PC3DOWNTO2_shadow_intermed_4 <= V_D_PC3DOWNTO2_shadow_intermed_3;
		V_D_PC3DOWNTO2_shadow_intermed_5 <= V_D_PC3DOWNTO2_shadow_intermed_4;
		RIN_D_PC3DOWNTO2_intermed_1 <= RIN.D.PC( 3 DOWNTO 2 );
		RIN_D_PC3DOWNTO2_intermed_2 <= RIN_D_PC3DOWNTO2_intermed_1;
		RIN_D_PC3DOWNTO2_intermed_3 <= RIN_D_PC3DOWNTO2_intermed_2;
		RIN_D_PC3DOWNTO2_intermed_4 <= RIN_D_PC3DOWNTO2_intermed_3;
		RIN_D_PC3DOWNTO2_intermed_5 <= RIN_D_PC3DOWNTO2_intermed_4;
		R_M_CTRL_PC3DOWNTO2_intermed_1 <= R.M.CTRL.PC( 3 DOWNTO 2 );
		R_E_CTRL_PC3DOWNTO2_intermed_1 <= R.E.CTRL.PC( 3 DOWNTO 2 );
		R_E_CTRL_PC3DOWNTO2_intermed_2 <= R_E_CTRL_PC3DOWNTO2_intermed_1;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC3DOWNTO2_shadow;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC3DOWNTO2_shadow_intermed_1;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_3 <= V_E_CTRL_PC3DOWNTO2_shadow_intermed_2;
		RIN_X_CTRL_PC3DOWNTO2_intermed_1 <= RIN.X.CTRL.PC( 3 DOWNTO 2 );
		R_A_CTRL_PC3DOWNTO2_intermed_1 <= R.A.CTRL.PC( 3 DOWNTO 2 );
		R_A_CTRL_PC3DOWNTO2_intermed_2 <= R_A_CTRL_PC3DOWNTO2_intermed_1;
		R_A_CTRL_PC3DOWNTO2_intermed_3 <= R_A_CTRL_PC3DOWNTO2_intermed_2;
		RIN_M_CTRL_PC3DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 3 DOWNTO 2 );
		RIN_M_CTRL_PC3DOWNTO2_intermed_2 <= RIN_M_CTRL_PC3DOWNTO2_intermed_1;
		RIN_A_CTRL_PC3DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 3 DOWNTO 2 );
		RIN_A_CTRL_PC3DOWNTO2_intermed_2 <= RIN_A_CTRL_PC3DOWNTO2_intermed_1;
		RIN_A_CTRL_PC3DOWNTO2_intermed_3 <= RIN_A_CTRL_PC3DOWNTO2_intermed_2;
		RIN_A_CTRL_PC3DOWNTO2_intermed_4 <= RIN_A_CTRL_PC3DOWNTO2_intermed_3;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC3DOWNTO2_shadow;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_2;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_4 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_3;
		V_M_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_M_CTRL_PC3DOWNTO2_shadow;
		V_M_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_M_CTRL_PC3DOWNTO2_shadow_intermed_1;
		RIN_E_CTRL_PC3DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 3 DOWNTO 2 );
		RIN_E_CTRL_PC3DOWNTO2_intermed_2 <= RIN_E_CTRL_PC3DOWNTO2_intermed_1;
		RIN_E_CTRL_PC3DOWNTO2_intermed_3 <= RIN_E_CTRL_PC3DOWNTO2_intermed_2;
		RIN_E_CTRL_RD6DOWNTO0_intermed_1 <= RIN.E.CTRL.RD( 6 DOWNTO 0 );
		RIN_E_CTRL_RD6DOWNTO0_intermed_2 <= RIN_E_CTRL_RD6DOWNTO0_intermed_1;
		RIN_M_CTRL_RD6DOWNTO0_intermed_1 <= RIN.M.CTRL.RD( 6 DOWNTO 0 );
		R_E_CTRL_RD6DOWNTO0_intermed_1 <= R.E.CTRL.RD( 6 DOWNTO 0 );
		V_E_CTRL_RD6DOWNTO0_shadow_intermed_1 <= V_E_CTRL_RD6DOWNTO0_shadow;
		V_E_CTRL_RD6DOWNTO0_shadow_intermed_2 <= V_E_CTRL_RD6DOWNTO0_shadow_intermed_1;
		V_A_CTRL_RD6DOWNTO0_shadow_intermed_1 <= V_A_CTRL_RD6DOWNTO0_shadow;
		V_A_CTRL_RD6DOWNTO0_shadow_intermed_2 <= V_A_CTRL_RD6DOWNTO0_shadow_intermed_1;
		V_A_CTRL_RD6DOWNTO0_shadow_intermed_3 <= V_A_CTRL_RD6DOWNTO0_shadow_intermed_2;
		R_A_CTRL_RD6DOWNTO0_intermed_1 <= R.A.CTRL.RD( 6 DOWNTO 0 );
		R_A_CTRL_RD6DOWNTO0_intermed_2 <= R_A_CTRL_RD6DOWNTO0_intermed_1;
		RIN_A_CTRL_RD6DOWNTO0_intermed_1 <= RIN.A.CTRL.RD( 6 DOWNTO 0 );
		RIN_A_CTRL_RD6DOWNTO0_intermed_2 <= RIN_A_CTRL_RD6DOWNTO0_intermed_1;
		RIN_A_CTRL_RD6DOWNTO0_intermed_3 <= RIN_A_CTRL_RD6DOWNTO0_intermed_2;
		RIN_A_CTRL_TT_intermed_1 <= RIN.A.CTRL.TT;
		RIN_A_CTRL_TT_intermed_2 <= RIN_A_CTRL_TT_intermed_1;
		R_A_CTRL_TT_intermed_1 <= R.A.CTRL.TT;
		RIN_E_CTRL_TT_intermed_1 <= RIN.E.CTRL.TT;
		V_A_CTRL_TT_shadow_intermed_1 <= V_A_CTRL_TT_shadow;
		V_A_CTRL_TT_shadow_intermed_2 <= V_A_CTRL_TT_shadow_intermed_1;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow;
		V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2 <= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1;
		R_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= R.X.RESULT( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= RIN.X.RESULT( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2 <= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1;
		RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1 <= RIN.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 );
		R_M_CTRL_TT3DOWNTO0_intermed_1 <= R.M.CTRL.TT( 3 DOWNTO 0 );
		R_A_CTRL_TT3DOWNTO0_intermed_1 <= R.A.CTRL.TT( 3 DOWNTO 0 );
		R_A_CTRL_TT3DOWNTO0_intermed_2 <= R_A_CTRL_TT3DOWNTO0_intermed_1;
		R_A_CTRL_TT3DOWNTO0_intermed_3 <= R_A_CTRL_TT3DOWNTO0_intermed_2;
		RIN_A_CTRL_TT3DOWNTO0_intermed_1 <= RIN.A.CTRL.TT( 3 DOWNTO 0 );
		RIN_A_CTRL_TT3DOWNTO0_intermed_2 <= RIN_A_CTRL_TT3DOWNTO0_intermed_1;
		RIN_A_CTRL_TT3DOWNTO0_intermed_3 <= RIN_A_CTRL_TT3DOWNTO0_intermed_2;
		RIN_A_CTRL_TT3DOWNTO0_intermed_4 <= RIN_A_CTRL_TT3DOWNTO0_intermed_3;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_A_CTRL_TT3DOWNTO0_shadow;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_1;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_3 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_2;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_4 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_3;
		R_E_CTRL_TT3DOWNTO0_intermed_1 <= R.E.CTRL.TT( 3 DOWNTO 0 );
		R_E_CTRL_TT3DOWNTO0_intermed_2 <= R_E_CTRL_TT3DOWNTO0_intermed_1;
		RIN_M_CTRL_TT3DOWNTO0_intermed_1 <= RIN.M.CTRL.TT( 3 DOWNTO 0 );
		RIN_M_CTRL_TT3DOWNTO0_intermed_2 <= RIN_M_CTRL_TT3DOWNTO0_intermed_1;
		V_M_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_M_CTRL_TT3DOWNTO0_shadow;
		V_M_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_M_CTRL_TT3DOWNTO0_shadow_intermed_1;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_E_CTRL_TT3DOWNTO0_shadow;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_E_CTRL_TT3DOWNTO0_shadow_intermed_1;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_3 <= V_E_CTRL_TT3DOWNTO0_shadow_intermed_2;
		RIN_X_CTRL_TT3DOWNTO0_intermed_1 <= RIN.X.CTRL.TT( 3 DOWNTO 0 );
		RIN_E_CTRL_TT3DOWNTO0_intermed_1 <= RIN.E.CTRL.TT( 3 DOWNTO 0 );
		RIN_E_CTRL_TT3DOWNTO0_intermed_2 <= RIN_E_CTRL_TT3DOWNTO0_intermed_1;
		RIN_E_CTRL_TT3DOWNTO0_intermed_3 <= RIN_E_CTRL_TT3DOWNTO0_intermed_2;
		R_M_CTRL_PC31DOWNTO12_intermed_1 <= R.M.CTRL.PC( 31 DOWNTO 12 );
		V_D_PC31DOWNTO12_shadow_intermed_1 <= V_D_PC31DOWNTO12_shadow;
		V_D_PC31DOWNTO12_shadow_intermed_2 <= V_D_PC31DOWNTO12_shadow_intermed_1;
		V_D_PC31DOWNTO12_shadow_intermed_3 <= V_D_PC31DOWNTO12_shadow_intermed_2;
		V_D_PC31DOWNTO12_shadow_intermed_4 <= V_D_PC31DOWNTO12_shadow_intermed_3;
		V_D_PC31DOWNTO12_shadow_intermed_5 <= V_D_PC31DOWNTO12_shadow_intermed_4;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO12_shadow;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_4 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_3;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO12_shadow;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_2;
		R_A_CTRL_PC31DOWNTO12_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 12 );
		R_A_CTRL_PC31DOWNTO12_intermed_2 <= R_A_CTRL_PC31DOWNTO12_intermed_1;
		R_A_CTRL_PC31DOWNTO12_intermed_3 <= R_A_CTRL_PC31DOWNTO12_intermed_2;
		R_E_CTRL_PC31DOWNTO12_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 12 );
		R_E_CTRL_PC31DOWNTO12_intermed_2 <= R_E_CTRL_PC31DOWNTO12_intermed_1;
		RIN_A_CTRL_PC31DOWNTO12_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 12 );
		RIN_A_CTRL_PC31DOWNTO12_intermed_2 <= RIN_A_CTRL_PC31DOWNTO12_intermed_1;
		RIN_A_CTRL_PC31DOWNTO12_intermed_3 <= RIN_A_CTRL_PC31DOWNTO12_intermed_2;
		RIN_A_CTRL_PC31DOWNTO12_intermed_4 <= RIN_A_CTRL_PC31DOWNTO12_intermed_3;
		RIN_E_CTRL_PC31DOWNTO12_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 12 );
		RIN_E_CTRL_PC31DOWNTO12_intermed_2 <= RIN_E_CTRL_PC31DOWNTO12_intermed_1;
		RIN_E_CTRL_PC31DOWNTO12_intermed_3 <= RIN_E_CTRL_PC31DOWNTO12_intermed_2;
		RIN_M_CTRL_PC31DOWNTO12_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 12 );
		RIN_M_CTRL_PC31DOWNTO12_intermed_2 <= RIN_M_CTRL_PC31DOWNTO12_intermed_1;
		R_D_PC31DOWNTO12_intermed_1 <= R.D.PC( 31 DOWNTO 12 );
		R_D_PC31DOWNTO12_intermed_2 <= R_D_PC31DOWNTO12_intermed_1;
		R_D_PC31DOWNTO12_intermed_3 <= R_D_PC31DOWNTO12_intermed_2;
		R_D_PC31DOWNTO12_intermed_4 <= R_D_PC31DOWNTO12_intermed_3;
		RIN_X_CTRL_PC31DOWNTO12_intermed_1 <= RIN.X.CTRL.PC( 31 DOWNTO 12 );
		RIN_D_PC31DOWNTO12_intermed_1 <= RIN.D.PC( 31 DOWNTO 12 );
		RIN_D_PC31DOWNTO12_intermed_2 <= RIN_D_PC31DOWNTO12_intermed_1;
		RIN_D_PC31DOWNTO12_intermed_3 <= RIN_D_PC31DOWNTO12_intermed_2;
		RIN_D_PC31DOWNTO12_intermed_4 <= RIN_D_PC31DOWNTO12_intermed_3;
		RIN_D_PC31DOWNTO12_intermed_5 <= RIN_D_PC31DOWNTO12_intermed_4;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_M_CTRL_PC31DOWNTO12_shadow;
		V_M_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_M_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_A_CTRL_RD7DOWNTO0_shadow_intermed_1 <= V_A_CTRL_RD7DOWNTO0_shadow;
		V_A_CTRL_RD7DOWNTO0_shadow_intermed_2 <= V_A_CTRL_RD7DOWNTO0_shadow_intermed_1;
		RIN_A_CTRL_RD7DOWNTO0_intermed_1 <= RIN.A.CTRL.RD ( 7 DOWNTO 0 );
		RIN_A_CTRL_RD7DOWNTO0_intermed_2 <= RIN_A_CTRL_RD7DOWNTO0_intermed_1;
		R_A_CTRL_RD7DOWNTO0_intermed_1 <= R.A.CTRL.RD ( 7 DOWNTO 0 );
		RIN_E_CTRL_RD7DOWNTO0_intermed_1 <= RIN.E.CTRL.RD ( 7 DOWNTO 0 );
		RIN_D_PC_intermed_1 <= RIN.D.PC;
		RIN_D_PC_intermed_2 <= RIN_D_PC_intermed_1;
		RIN_D_PC_intermed_3 <= RIN_D_PC_intermed_2;
		RIN_A_CTRL_PC_intermed_1 <= RIN.A.CTRL.PC;
		RIN_A_CTRL_PC_intermed_2 <= RIN_A_CTRL_PC_intermed_1;
		R_A_CTRL_PC_intermed_1 <= R.A.CTRL.PC;
		V_A_CTRL_PC_shadow_intermed_1 <= V_A_CTRL_PC_shadow;
		V_A_CTRL_PC_shadow_intermed_2 <= V_A_CTRL_PC_shadow_intermed_1;
		R_D_PC_intermed_1 <= R.D.PC;
		R_D_PC_intermed_2 <= R_D_PC_intermed_1;
		RIN_E_CTRL_PC_intermed_1 <= RIN.E.CTRL.PC;
		V_D_PC_shadow_intermed_1 <= V_D_PC_shadow;
		V_D_PC_shadow_intermed_2 <= V_D_PC_shadow_intermed_1;
		V_D_PC_shadow_intermed_3 <= V_D_PC_shadow_intermed_2;
		V_D_PC31DOWNTO2_shadow_intermed_1 <= V_D_PC31DOWNTO2_shadow;
		V_D_PC31DOWNTO2_shadow_intermed_2 <= V_D_PC31DOWNTO2_shadow_intermed_1;
		V_D_PC31DOWNTO2_shadow_intermed_3 <= V_D_PC31DOWNTO2_shadow_intermed_2;
		RIN_D_PC31DOWNTO2_intermed_1 <= RIN.D.PC( 31 DOWNTO 2 );
		RIN_D_PC31DOWNTO2_intermed_2 <= RIN_D_PC31DOWNTO2_intermed_1;
		RIN_D_PC31DOWNTO2_intermed_3 <= RIN_D_PC31DOWNTO2_intermed_2;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO2_shadow;
		V_A_CTRL_PC31DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1;
		R_D_PC31DOWNTO2_intermed_1 <= R.D.PC( 31 DOWNTO 2 );
		R_D_PC31DOWNTO2_intermed_2 <= R_D_PC31DOWNTO2_intermed_1;
		RIN_A_CTRL_PC31DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO2_intermed_2 <= RIN_A_CTRL_PC31DOWNTO2_intermed_1;
		R_A_CTRL_PC31DOWNTO2_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 2 );
		RIN_E_CTRL_PC31DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 2 );
		RIN_A_CTRL_PC31DOWNTO4_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 4 );
		RIN_A_CTRL_PC31DOWNTO4_intermed_2 <= RIN_A_CTRL_PC31DOWNTO4_intermed_1;
		RIN_A_CTRL_PC31DOWNTO4_intermed_3 <= RIN_A_CTRL_PC31DOWNTO4_intermed_2;
		R_A_CTRL_PC31DOWNTO4_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 4 );
		R_A_CTRL_PC31DOWNTO4_intermed_2 <= R_A_CTRL_PC31DOWNTO4_intermed_1;
		R_D_PC31DOWNTO4_intermed_1 <= R.D.PC( 31 DOWNTO 4 );
		R_D_PC31DOWNTO4_intermed_2 <= R_D_PC31DOWNTO4_intermed_1;
		R_D_PC31DOWNTO4_intermed_3 <= R_D_PC31DOWNTO4_intermed_2;
		V_D_PC31DOWNTO4_shadow_intermed_1 <= V_D_PC31DOWNTO4_shadow;
		V_D_PC31DOWNTO4_shadow_intermed_2 <= V_D_PC31DOWNTO4_shadow_intermed_1;
		V_D_PC31DOWNTO4_shadow_intermed_3 <= V_D_PC31DOWNTO4_shadow_intermed_2;
		V_D_PC31DOWNTO4_shadow_intermed_4 <= V_D_PC31DOWNTO4_shadow_intermed_3;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO4_shadow;
		V_E_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO4_shadow_intermed_1;
		RIN_M_CTRL_PC31DOWNTO4_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 4 );
		RIN_D_PC31DOWNTO4_intermed_1 <= RIN.D.PC( 31 DOWNTO 4 );
		RIN_D_PC31DOWNTO4_intermed_2 <= RIN_D_PC31DOWNTO4_intermed_1;
		RIN_D_PC31DOWNTO4_intermed_3 <= RIN_D_PC31DOWNTO4_intermed_2;
		RIN_D_PC31DOWNTO4_intermed_4 <= RIN_D_PC31DOWNTO4_intermed_3;
		RIN_E_CTRL_PC31DOWNTO4_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 4 );
		RIN_E_CTRL_PC31DOWNTO4_intermed_2 <= RIN_E_CTRL_PC31DOWNTO4_intermed_1;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO4_shadow;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_2;
		R_E_CTRL_PC31DOWNTO4_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 4 );
		R_D_PC3DOWNTO2_intermed_1 <= R.D.PC( 3 DOWNTO 2 );
		R_D_PC3DOWNTO2_intermed_2 <= R_D_PC3DOWNTO2_intermed_1;
		R_D_PC3DOWNTO2_intermed_3 <= R_D_PC3DOWNTO2_intermed_2;
		V_D_PC3DOWNTO2_shadow_intermed_1 <= V_D_PC3DOWNTO2_shadow;
		V_D_PC3DOWNTO2_shadow_intermed_2 <= V_D_PC3DOWNTO2_shadow_intermed_1;
		V_D_PC3DOWNTO2_shadow_intermed_3 <= V_D_PC3DOWNTO2_shadow_intermed_2;
		V_D_PC3DOWNTO2_shadow_intermed_4 <= V_D_PC3DOWNTO2_shadow_intermed_3;
		RIN_D_PC3DOWNTO2_intermed_1 <= RIN.D.PC( 3 DOWNTO 2 );
		RIN_D_PC3DOWNTO2_intermed_2 <= RIN_D_PC3DOWNTO2_intermed_1;
		RIN_D_PC3DOWNTO2_intermed_3 <= RIN_D_PC3DOWNTO2_intermed_2;
		RIN_D_PC3DOWNTO2_intermed_4 <= RIN_D_PC3DOWNTO2_intermed_3;
		R_E_CTRL_PC3DOWNTO2_intermed_1 <= R.E.CTRL.PC( 3 DOWNTO 2 );
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_E_CTRL_PC3DOWNTO2_shadow;
		V_E_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_E_CTRL_PC3DOWNTO2_shadow_intermed_1;
		R_A_CTRL_PC3DOWNTO2_intermed_1 <= R.A.CTRL.PC( 3 DOWNTO 2 );
		R_A_CTRL_PC3DOWNTO2_intermed_2 <= R_A_CTRL_PC3DOWNTO2_intermed_1;
		RIN_M_CTRL_PC3DOWNTO2_intermed_1 <= RIN.M.CTRL.PC( 3 DOWNTO 2 );
		RIN_A_CTRL_PC3DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 3 DOWNTO 2 );
		RIN_A_CTRL_PC3DOWNTO2_intermed_2 <= RIN_A_CTRL_PC3DOWNTO2_intermed_1;
		RIN_A_CTRL_PC3DOWNTO2_intermed_3 <= RIN_A_CTRL_PC3DOWNTO2_intermed_2;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC3DOWNTO2_shadow;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_1;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_3 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_2;
		RIN_E_CTRL_PC3DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 3 DOWNTO 2 );
		RIN_E_CTRL_PC3DOWNTO2_intermed_2 <= RIN_E_CTRL_PC3DOWNTO2_intermed_1;
		RIN_E_CTRL_RD6DOWNTO0_intermed_1 <= RIN.E.CTRL.RD( 6 DOWNTO 0 );
		V_A_CTRL_RD6DOWNTO0_shadow_intermed_1 <= V_A_CTRL_RD6DOWNTO0_shadow;
		V_A_CTRL_RD6DOWNTO0_shadow_intermed_2 <= V_A_CTRL_RD6DOWNTO0_shadow_intermed_1;
		R_A_CTRL_RD6DOWNTO0_intermed_1 <= R.A.CTRL.RD( 6 DOWNTO 0 );
		RIN_A_CTRL_RD6DOWNTO0_intermed_1 <= RIN.A.CTRL.RD( 6 DOWNTO 0 );
		RIN_A_CTRL_RD6DOWNTO0_intermed_2 <= RIN_A_CTRL_RD6DOWNTO0_intermed_1;
		R_A_CTRL_TT3DOWNTO0_intermed_1 <= R.A.CTRL.TT( 3 DOWNTO 0 );
		R_A_CTRL_TT3DOWNTO0_intermed_2 <= R_A_CTRL_TT3DOWNTO0_intermed_1;
		RIN_A_CTRL_TT3DOWNTO0_intermed_1 <= RIN.A.CTRL.TT( 3 DOWNTO 0 );
		RIN_A_CTRL_TT3DOWNTO0_intermed_2 <= RIN_A_CTRL_TT3DOWNTO0_intermed_1;
		RIN_A_CTRL_TT3DOWNTO0_intermed_3 <= RIN_A_CTRL_TT3DOWNTO0_intermed_2;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_A_CTRL_TT3DOWNTO0_shadow;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_1;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_3 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_2;
		R_E_CTRL_TT3DOWNTO0_intermed_1 <= R.E.CTRL.TT( 3 DOWNTO 0 );
		RIN_M_CTRL_TT3DOWNTO0_intermed_1 <= RIN.M.CTRL.TT( 3 DOWNTO 0 );
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_E_CTRL_TT3DOWNTO0_shadow;
		V_E_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_E_CTRL_TT3DOWNTO0_shadow_intermed_1;
		RIN_E_CTRL_TT3DOWNTO0_intermed_1 <= RIN.E.CTRL.TT( 3 DOWNTO 0 );
		RIN_E_CTRL_TT3DOWNTO0_intermed_2 <= RIN_E_CTRL_TT3DOWNTO0_intermed_1;
		V_D_PC31DOWNTO12_shadow_intermed_1 <= V_D_PC31DOWNTO12_shadow;
		V_D_PC31DOWNTO12_shadow_intermed_2 <= V_D_PC31DOWNTO12_shadow_intermed_1;
		V_D_PC31DOWNTO12_shadow_intermed_3 <= V_D_PC31DOWNTO12_shadow_intermed_2;
		V_D_PC31DOWNTO12_shadow_intermed_4 <= V_D_PC31DOWNTO12_shadow_intermed_3;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO12_shadow;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_1;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_3 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_2;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_E_CTRL_PC31DOWNTO12_shadow;
		V_E_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_E_CTRL_PC31DOWNTO12_shadow_intermed_1;
		R_A_CTRL_PC31DOWNTO12_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 12 );
		R_A_CTRL_PC31DOWNTO12_intermed_2 <= R_A_CTRL_PC31DOWNTO12_intermed_1;
		R_E_CTRL_PC31DOWNTO12_intermed_1 <= R.E.CTRL.PC( 31 DOWNTO 12 );
		RIN_A_CTRL_PC31DOWNTO12_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 12 );
		RIN_A_CTRL_PC31DOWNTO12_intermed_2 <= RIN_A_CTRL_PC31DOWNTO12_intermed_1;
		RIN_A_CTRL_PC31DOWNTO12_intermed_3 <= RIN_A_CTRL_PC31DOWNTO12_intermed_2;
		RIN_E_CTRL_PC31DOWNTO12_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 12 );
		RIN_E_CTRL_PC31DOWNTO12_intermed_2 <= RIN_E_CTRL_PC31DOWNTO12_intermed_1;
		RIN_M_CTRL_PC31DOWNTO12_intermed_1 <= RIN.M.CTRL.PC( 31 DOWNTO 12 );
		R_D_PC31DOWNTO12_intermed_1 <= R.D.PC( 31 DOWNTO 12 );
		R_D_PC31DOWNTO12_intermed_2 <= R_D_PC31DOWNTO12_intermed_1;
		R_D_PC31DOWNTO12_intermed_3 <= R_D_PC31DOWNTO12_intermed_2;
		RIN_D_PC31DOWNTO12_intermed_1 <= RIN.D.PC( 31 DOWNTO 12 );
		RIN_D_PC31DOWNTO12_intermed_2 <= RIN_D_PC31DOWNTO12_intermed_1;
		RIN_D_PC31DOWNTO12_intermed_3 <= RIN_D_PC31DOWNTO12_intermed_2;
		RIN_D_PC31DOWNTO12_intermed_4 <= RIN_D_PC31DOWNTO12_intermed_3;
		RIN_A_CTRL_PC31DOWNTO4_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 4 );
		RIN_A_CTRL_PC31DOWNTO4_intermed_2 <= RIN_A_CTRL_PC31DOWNTO4_intermed_1;
		R_A_CTRL_PC31DOWNTO4_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 4 );
		R_D_PC31DOWNTO4_intermed_1 <= R.D.PC( 31 DOWNTO 4 );
		R_D_PC31DOWNTO4_intermed_2 <= R_D_PC31DOWNTO4_intermed_1;
		V_D_PC31DOWNTO4_shadow_intermed_1 <= V_D_PC31DOWNTO4_shadow;
		V_D_PC31DOWNTO4_shadow_intermed_2 <= V_D_PC31DOWNTO4_shadow_intermed_1;
		V_D_PC31DOWNTO4_shadow_intermed_3 <= V_D_PC31DOWNTO4_shadow_intermed_2;
		RIN_D_PC31DOWNTO4_intermed_1 <= RIN.D.PC( 31 DOWNTO 4 );
		RIN_D_PC31DOWNTO4_intermed_2 <= RIN_D_PC31DOWNTO4_intermed_1;
		RIN_D_PC31DOWNTO4_intermed_3 <= RIN_D_PC31DOWNTO4_intermed_2;
		RIN_E_CTRL_PC31DOWNTO4_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 4 );
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO4_shadow;
		V_A_CTRL_PC31DOWNTO4_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO4_shadow_intermed_1;
		R_D_PC3DOWNTO2_intermed_1 <= R.D.PC( 3 DOWNTO 2 );
		R_D_PC3DOWNTO2_intermed_2 <= R_D_PC3DOWNTO2_intermed_1;
		V_D_PC3DOWNTO2_shadow_intermed_1 <= V_D_PC3DOWNTO2_shadow;
		V_D_PC3DOWNTO2_shadow_intermed_2 <= V_D_PC3DOWNTO2_shadow_intermed_1;
		V_D_PC3DOWNTO2_shadow_intermed_3 <= V_D_PC3DOWNTO2_shadow_intermed_2;
		RIN_D_PC3DOWNTO2_intermed_1 <= RIN.D.PC( 3 DOWNTO 2 );
		RIN_D_PC3DOWNTO2_intermed_2 <= RIN_D_PC3DOWNTO2_intermed_1;
		RIN_D_PC3DOWNTO2_intermed_3 <= RIN_D_PC3DOWNTO2_intermed_2;
		R_A_CTRL_PC3DOWNTO2_intermed_1 <= R.A.CTRL.PC( 3 DOWNTO 2 );
		RIN_A_CTRL_PC3DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 3 DOWNTO 2 );
		RIN_A_CTRL_PC3DOWNTO2_intermed_2 <= RIN_A_CTRL_PC3DOWNTO2_intermed_1;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_1 <= V_A_CTRL_PC3DOWNTO2_shadow;
		V_A_CTRL_PC3DOWNTO2_shadow_intermed_2 <= V_A_CTRL_PC3DOWNTO2_shadow_intermed_1;
		RIN_E_CTRL_PC3DOWNTO2_intermed_1 <= RIN.E.CTRL.PC( 3 DOWNTO 2 );
		R_A_CTRL_TT3DOWNTO0_intermed_1 <= R.A.CTRL.TT( 3 DOWNTO 0 );
		RIN_A_CTRL_TT3DOWNTO0_intermed_1 <= RIN.A.CTRL.TT( 3 DOWNTO 0 );
		RIN_A_CTRL_TT3DOWNTO0_intermed_2 <= RIN_A_CTRL_TT3DOWNTO0_intermed_1;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_1 <= V_A_CTRL_TT3DOWNTO0_shadow;
		V_A_CTRL_TT3DOWNTO0_shadow_intermed_2 <= V_A_CTRL_TT3DOWNTO0_shadow_intermed_1;
		RIN_E_CTRL_TT3DOWNTO0_intermed_1 <= RIN.E.CTRL.TT( 3 DOWNTO 0 );
		V_D_PC31DOWNTO12_shadow_intermed_1 <= V_D_PC31DOWNTO12_shadow;
		V_D_PC31DOWNTO12_shadow_intermed_2 <= V_D_PC31DOWNTO12_shadow_intermed_1;
		V_D_PC31DOWNTO12_shadow_intermed_3 <= V_D_PC31DOWNTO12_shadow_intermed_2;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_1 <= V_A_CTRL_PC31DOWNTO12_shadow;
		V_A_CTRL_PC31DOWNTO12_shadow_intermed_2 <= V_A_CTRL_PC31DOWNTO12_shadow_intermed_1;
		R_A_CTRL_PC31DOWNTO12_intermed_1 <= R.A.CTRL.PC( 31 DOWNTO 12 );
		RIN_A_CTRL_PC31DOWNTO12_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 12 );
		RIN_A_CTRL_PC31DOWNTO12_intermed_2 <= RIN_A_CTRL_PC31DOWNTO12_intermed_1;
		RIN_E_CTRL_PC31DOWNTO12_intermed_1 <= RIN.E.CTRL.PC( 31 DOWNTO 12 );
		R_D_PC31DOWNTO12_intermed_1 <= R.D.PC( 31 DOWNTO 12 );
		R_D_PC31DOWNTO12_intermed_2 <= R_D_PC31DOWNTO12_intermed_1;
		RIN_D_PC31DOWNTO12_intermed_1 <= RIN.D.PC( 31 DOWNTO 12 );
		RIN_D_PC31DOWNTO12_intermed_2 <= RIN_D_PC31DOWNTO12_intermed_1;
		RIN_D_PC31DOWNTO12_intermed_3 <= RIN_D_PC31DOWNTO12_intermed_2;
		RIN_A_CTRL_PC31DOWNTO4_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 4 );
		R_D_PC31DOWNTO4_intermed_1 <= R.D.PC( 31 DOWNTO 4 );
		V_D_PC31DOWNTO4_shadow_intermed_1 <= V_D_PC31DOWNTO4_shadow;
		V_D_PC31DOWNTO4_shadow_intermed_2 <= V_D_PC31DOWNTO4_shadow_intermed_1;
		RIN_D_PC31DOWNTO4_intermed_1 <= RIN.D.PC( 31 DOWNTO 4 );
		RIN_D_PC31DOWNTO4_intermed_2 <= RIN_D_PC31DOWNTO4_intermed_1;
		R_D_PC3DOWNTO2_intermed_1 <= R.D.PC( 3 DOWNTO 2 );
		V_D_PC3DOWNTO2_shadow_intermed_1 <= V_D_PC3DOWNTO2_shadow;
		V_D_PC3DOWNTO2_shadow_intermed_2 <= V_D_PC3DOWNTO2_shadow_intermed_1;
		RIN_D_PC3DOWNTO2_intermed_1 <= RIN.D.PC( 3 DOWNTO 2 );
		RIN_D_PC3DOWNTO2_intermed_2 <= RIN_D_PC3DOWNTO2_intermed_1;
		RIN_A_CTRL_PC3DOWNTO2_intermed_1 <= RIN.A.CTRL.PC( 3 DOWNTO 2 );
		V_D_PC31DOWNTO12_shadow_intermed_1 <= V_D_PC31DOWNTO12_shadow;
		V_D_PC31DOWNTO12_shadow_intermed_2 <= V_D_PC31DOWNTO12_shadow_intermed_1;
		RIN_A_CTRL_PC31DOWNTO12_intermed_1 <= RIN.A.CTRL.PC( 31 DOWNTO 12 );
		R_D_PC31DOWNTO12_intermed_1 <= R.D.PC( 31 DOWNTO 12 );
		RIN_D_PC31DOWNTO12_intermed_1 <= RIN.D.PC( 31 DOWNTO 12 );
		RIN_D_PC31DOWNTO12_intermed_2 <= RIN_D_PC31DOWNTO12_intermed_1;
	end if;
end process;

dfp_trap_vector(0) <= '1' when (RP.ERROR /= '1') else '0';
dfp_trap_vector(1) <= '1' when (RP.ERROR /= '0') else '0';
dfp_trap_vector(2) <= '1' when (RP.ERROR /= RPIN_ERROR_intermed_1) else '0';
dfp_trap_vector(3) <= '1' when (RP.ERROR /= VP_ERROR_shadow_intermed_1) else '0';
dfp_trap_vector(4) <= '1' when (R.W.S.S /= V_W_S_S_shadow_intermed_1) else '0';
dfp_trap_vector(5) <= '1' when (R.W.S.S /= '1') else '0';
dfp_trap_vector(6) <= '1' when (R.W.S.S /= RIN_W_S_S_intermed_1) else '0';
dfp_trap_vector(7) <= '1' when (R.W.S.PS /= V_W_S_S_shadow_intermed_2) else '0';
dfp_trap_vector(8) <= '1' when (R.W.S.PS /= V_W_S_PS_shadow_intermed_1) else '0';
dfp_trap_vector(9) <= '1' when (R.W.S.PS /= '1') else '0';
dfp_trap_vector(10) <= '1' when (R.W.S.PS /= RIN_W_S_PS_intermed_1) else '0';
dfp_trap_vector(11) <= '1' when (R.W.S.PS /= R_W_S_S_intermed_1) else '0';
dfp_trap_vector(12) <= '1' when (R.W.S.PS /= RIN_W_S_S_intermed_2) else '0';
dfp_trap_vector(13) <= '1' when (R.X.RESULT ( 6 DOWNTO 0 ) /= R_X_RESULT6DOWNTO0_intermed_2) else '0';
dfp_trap_vector(14) <= '1' when (R.X.RESULT ( 6 DOWNTO 0 ) /= V_X_RESULT6DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(15) <= '1' when (R.X.RESULT ( 6 DOWNTO 0 ) /= V_X_RESULT6DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(16) <= '1' when (R.X.RESULT ( 6 DOWNTO 0 ) /= RIN_X_RESULT6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(17) <= '1' when (R.X.RESULT ( 6 DOWNTO 0 ) /= RIN_X_RESULT6DOWNTO0_intermed_2) else '0';
dfp_trap_vector(18) <= '1' when (R.X.DATA ( 0 ) /= V_X_DATA0_shadow_intermed_2) else '0';
dfp_trap_vector(19) <= '1' when (R.X.DATA ( 0 ) /= R_X_DATA0_intermed_2) else '0';
dfp_trap_vector(20) <= '1' when (R.X.DATA ( 0 ) /= DCO_DATA0_intermed_1) else '0';
dfp_trap_vector(21) <= '1' when (R.X.DATA ( 0 ) /= V_X_DATA0_shadow_intermed_1) else '0';
dfp_trap_vector(22) <= '1' when (R.X.DATA ( 0 ) /= RIN_X_DATA0_intermed_1) else '0';
dfp_trap_vector(23) <= '1' when (R.X.DATA ( 0 ) /= RIN_X_DATA0_intermed_2) else '0';
dfp_trap_vector(24) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= R_M_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(25) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_M_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(26) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(27) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_A_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(28) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= V_X_CTRL_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(29) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(30) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= R_A_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(31) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(32) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= R_A_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(33) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= R_X_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(34) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= R_E_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(35) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= V_D_PC31DOWNTO2_shadow_intermed_6) else '0';
dfp_trap_vector(36) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_D_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(37) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_E_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(38) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_A_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(39) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_X_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(40) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_X_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(41) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_M_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(42) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(43) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= R_E_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(44) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(45) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= R_D_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(46) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= R_M_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(47) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_E_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(48) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= V_X_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(49) <= '1' when (R.X.CTRL.PC ( 31 DOWNTO 2 ) /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(50) <= '1' when (RFI.WREN /= DCO.SCANEN) else '0';
dfp_trap_vector(51) <= '1' when (RFI.WREN /= V_X_ANNUL_ALL_shadow_intermed_4) else '0';
dfp_trap_vector(52) <= '1' when (RFI.WREN /= RIN_A_CTRL_ANNUL_intermed_5) else '0';
dfp_trap_vector(53) <= '1' when (RFI.WREN /= R_M_CTRL_WREG_intermed_1) else '0';
dfp_trap_vector(54) <= '1' when (RFI.WREN /= R.X.CTRL.WREG) else '0';
dfp_trap_vector(55) <= '1' when (RFI.WREN /= R_A_CTRL_ANNUL_intermed_4) else '0';
dfp_trap_vector(56) <= '1' when (RFI.WREN /= RIN_X_ANNUL_ALL_intermed_5) else '0';
dfp_trap_vector(57) <= '1' when (RFI.WREN /= V_M_CTRL_WREG_shadow_intermed_2) else '0';
dfp_trap_vector(58) <= '1' when (RFI.WREN /= R_X_ANNUL_ALL_intermed_4) else '0';
dfp_trap_vector(59) <= '1' when (RFI.WREN /= HOLDN) else '0';
dfp_trap_vector(60) <= '1' when (RFI.WREN /= V_X_CTRL_WREG_shadow_intermed_1) else '0';
dfp_trap_vector(61) <= '1' when (RFI.WREN /= R_E_CTRL_WREG_intermed_2) else '0';
dfp_trap_vector(62) <= '1' when (RFI.WREN /= RIN_X_CTRL_WREG_intermed_1) else '0';
dfp_trap_vector(63) <= '1' when (RFI.WREN /= '1') else '0';
dfp_trap_vector(64) <= '1' when (RFI.WREN /= '0') else '0';
dfp_trap_vector(65) <= '1' when (RFI.WREN /= XC_WREG_shadow) else '0';
dfp_trap_vector(66) <= '1' when (RFI.WREN /= V_A_CTRL_ANNUL_shadow_intermed_4) else '0';
dfp_trap_vector(67) <= '1' when (RFI.WREN /= RIN_E_CTRL_WREG_intermed_3) else '0';
dfp_trap_vector(68) <= '1' when (RFI.WREN /= RIN_M_CTRL_WREG_intermed_2) else '0';
dfp_trap_vector(69) <= '1' when (RFI.WREN /= V_E_CTRL_WREG_shadow_intermed_3) else '0';
dfp_trap_vector(70) <= '1' when (RFI.WREN /= RIN_A_CTRL_WREG_intermed_4) else '0';
dfp_trap_vector(71) <= '1' when (RFI.WREN /= V_A_CTRL_WREG_shadow_intermed_4) else '0';
dfp_trap_vector(72) <= '1' when (RFI.WREN /= R_A_CTRL_WREG_intermed_3) else '0';
dfp_trap_vector(73) <= '1' when (IRQO.INTACK /= RIN_X_INTACK_intermed_1) else '0';
dfp_trap_vector(74) <= '1' when (IRQO.INTACK /= V_X_INTACK_shadow_intermed_1) else '0';
dfp_trap_vector(75) <= '1' when (IRQO.INTACK /= HOLDN) else '0';
dfp_trap_vector(76) <= '1' when (IRQO.INTACK /= R.X.INTACK) else '0';
dfp_trap_vector(77) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= V_X_CTRL_TT3DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(78) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= R_M_CTRL_TT3DOWNTO0_intermed_3) else '0';
dfp_trap_vector(79) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= V_M_CTRL_TT3DOWNTO0_shadow_intermed_4) else '0';
dfp_trap_vector(80) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_4) else '0';
dfp_trap_vector(81) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= R_X_RESULT6DOWNTO03DOWNTO0_intermed_3) else '0';
dfp_trap_vector(82) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= R_A_CTRL_TT3DOWNTO0_intermed_5) else '0';
dfp_trap_vector(83) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= RIN_A_CTRL_TT3DOWNTO0_intermed_6) else '0';
dfp_trap_vector(84) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_4) else '0';
dfp_trap_vector(85) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= V_A_CTRL_TT3DOWNTO0_shadow_intermed_6) else '0';
dfp_trap_vector(86) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_3) else '0';
dfp_trap_vector(87) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= R_W_S_TT3DOWNTO0_intermed_2) else '0';
dfp_trap_vector(88) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= R_X_RESULT6DOWNTO03DOWNTO0_intermed_2) else '0';
dfp_trap_vector(89) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= R_E_CTRL_TT3DOWNTO0_intermed_4) else '0';
dfp_trap_vector(90) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(91) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= RIN_W_S_TT3DOWNTO0_intermed_2) else '0';
dfp_trap_vector(92) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= V_E_CTRL_TT3DOWNTO0_shadow_intermed_5) else '0';
dfp_trap_vector(93) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= RIN_W_S_TT3DOWNTO0_intermed_1) else '0';
dfp_trap_vector(94) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= RIN_M_CTRL_TT3DOWNTO0_intermed_4) else '0';
dfp_trap_vector(95) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= RIN_X_CTRL_TT3DOWNTO0_intermed_3) else '0';
dfp_trap_vector(96) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= V_W_S_TT3DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(97) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= R_X_CTRL_TT3DOWNTO0_intermed_2) else '0';
dfp_trap_vector(98) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= RIN_E_CTRL_TT3DOWNTO0_intermed_5) else '0';
dfp_trap_vector(99) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= V_W_S_TT3DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(100) <= '1' when (R.W.S.TT ( 3 DOWNTO 0 ) /= XC_VECTT3DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(101) <= '1' when (DCI.INTACK /= RIN_X_INTACK_intermed_1) else '0';
dfp_trap_vector(102) <= '1' when (DCI.INTACK /= V_X_INTACK_shadow_intermed_1) else '0';
dfp_trap_vector(103) <= '1' when (DCI.INTACK /= HOLDN) else '0';
dfp_trap_vector(104) <= '1' when (DCI.INTACK /= R.X.INTACK) else '0';
dfp_trap_vector(105) <= '1' when (R.M.RESULT ( 1 DOWNTO 0 ) /= V_M_RESULT1DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(106) <= '1' when (R.M.RESULT ( 1 DOWNTO 0 ) /= RIN_M_RESULT1DOWNTO0_intermed_1) else '0';
dfp_trap_vector(107) <= '1' when (R.M.RESULT ( 1 DOWNTO 0 ) /= RIN_M_RESULT1DOWNTO0_intermed_2) else '0';
dfp_trap_vector(108) <= '1' when (R.M.RESULT ( 1 DOWNTO 0 ) /= V_M_RESULT1DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(109) <= '1' when (R.M.RESULT ( 1 DOWNTO 0 ) /= R_M_RESULT1DOWNTO0_intermed_2) else '0';
dfp_trap_vector(110) <= '1' when (DCI.LOCK /= V_X_ANNUL_ALL_shadow_intermed_1) else '0';
dfp_trap_vector(111) <= '1' when (DCI.LOCK /= RIN_A_CTRL_ANNUL_intermed_3) else '0';
dfp_trap_vector(112) <= '1' when (DCI.LOCK /= RIN_E_CTRL_ANNUL_intermed_2) else '0';
dfp_trap_vector(113) <= '1' when (DCI.LOCK /= R_A_CTRL_ANNUL_intermed_2) else '0';
dfp_trap_vector(114) <= '1' when (DCI.LOCK /= V_M_CTRL_ANNUL_shadow_intermed_1) else '0';
dfp_trap_vector(115) <= '1' when (DCI.LOCK /= RIN_X_ANNUL_ALL_intermed_2) else '0';
dfp_trap_vector(116) <= '1' when (DCI.LOCK /= R_X_ANNUL_ALL_intermed_1) else '0';
dfp_trap_vector(117) <= '1' when (DCI.LOCK /= R.M.CTRL.ANNUL) else '0';
dfp_trap_vector(118) <= '1' when (DCI.LOCK /= RIN_M_DCI_LOCK_intermed_1) else '0';
dfp_trap_vector(119) <= '1' when (DCI.LOCK /= '1') else '0';
dfp_trap_vector(120) <= '1' when (DCI.LOCK /= V_E_CTRL_ANNUL_shadow_intermed_2) else '0';
dfp_trap_vector(121) <= '1' when (DCI.LOCK /= '0') else '0';
dfp_trap_vector(122) <= '1' when (DCI.LOCK /= V_A_CTRL_ANNUL_shadow_intermed_3) else '0';
dfp_trap_vector(123) <= '1' when (DCI.LOCK /= RIN_M_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(124) <= '1' when (DCI.LOCK /= R.M.DCI.LOCK) else '0';
dfp_trap_vector(125) <= '1' when (DCI.LOCK /= R_E_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(126) <= '1' when (DCI.LOCK /= V_M_DCI_LOCK_shadow_intermed_1) else '0';
dfp_trap_vector(127) <= '1' when (R.X.DATA ( 0 ) ( 31 ) /= RIN_X_DATA031_intermed_2) else '0';
dfp_trap_vector(128) <= '1' when (R.X.DATA ( 0 ) ( 31 ) /= V_X_DATA031_shadow_intermed_2) else '0';
dfp_trap_vector(129) <= '1' when (R.X.DATA ( 0 ) ( 31 ) /= V_X_DATA031_shadow_intermed_2) else '0';
dfp_trap_vector(130) <= '1' when (R.X.DATA ( 0 ) ( 31 ) /= RIN_X_DATA031_intermed_2) else '0';
dfp_trap_vector(131) <= '1' when (R.X.DATA ( 0 ) ( 31 ) /= RIN_X_DATA031_intermed_1) else '0';
dfp_trap_vector(132) <= '1' when (R.X.DATA ( 0 ) ( 31 ) /= DCO_DATA031_intermed_2) else '0';
dfp_trap_vector(133) <= '1' when (R.X.DATA ( 0 ) ( 31 ) /= R_X_DATA031_intermed_2) else '0';
dfp_trap_vector(134) <= '1' when (R.X.DATA ( 0 ) ( 31 ) /= R_X_DATA031_intermed_2) else '0';
dfp_trap_vector(135) <= '1' when (R.X.DATA ( 0 ) ( 31 ) /= V_X_DATA031_shadow_intermed_1) else '0';
dfp_trap_vector(136) <= '1' when (R.E.CTRL.INST ( 19 ) /= DE_INST19_shadow_intermed_3) else '0';
dfp_trap_vector(137) <= '1' when (R.E.CTRL.INST ( 19 ) /= V_A_CTRL_INST19_shadow_intermed_3) else '0';
dfp_trap_vector(138) <= '1' when (R.E.CTRL.INST ( 19 ) /= V_E_CTRL_INST19_shadow_intermed_1) else '0';
dfp_trap_vector(139) <= '1' when (R.E.CTRL.INST ( 19 ) /= V_E_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(140) <= '1' when (R.E.CTRL.INST ( 19 ) /= R_E_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(141) <= '1' when (R.E.CTRL.INST ( 19 ) /= RIN_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(142) <= '1' when (R.E.CTRL.INST ( 19 ) /= R_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(143) <= '1' when (R.E.CTRL.INST ( 19 ) /= R_A_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(144) <= '1' when (R.E.CTRL.INST ( 19 ) /= RIN_A_CTRL_INST19_intermed_3) else '0';
dfp_trap_vector(145) <= '1' when (R.E.CTRL.INST ( 19 ) /= RIN_E_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(146) <= '1' when (R.E.CTRL.INST ( 19 ) /= RIN_E_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(147) <= '1' when (R.E.CTRL.INST ( 19 ) /= V_A_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(148) <= '1' when (R.E.CTRL.INST ( 20 ) /= V_A_CTRL_INST20_shadow_intermed_2) else '0';
dfp_trap_vector(149) <= '1' when (R.E.CTRL.INST ( 20 ) /= RIN_A_CTRL_INST20_intermed_2) else '0';
dfp_trap_vector(150) <= '1' when (R.E.CTRL.INST ( 20 ) /= RIN_E_CTRL_INST20_intermed_1) else '0';
dfp_trap_vector(151) <= '1' when (R.E.CTRL.INST ( 20 ) /= R_A_CTRL_INST20_intermed_1) else '0';
dfp_trap_vector(152) <= '1' when (R.E.CTRL.INST ( 20 ) /= R_E_CTRL_INST20_intermed_2) else '0';
dfp_trap_vector(153) <= '1' when (R.E.CTRL.INST ( 20 ) /= RIN_A_CTRL_INST20_intermed_3) else '0';
dfp_trap_vector(154) <= '1' when (R.E.CTRL.INST ( 20 ) /= V_E_CTRL_INST20_shadow_intermed_2) else '0';
dfp_trap_vector(155) <= '1' when (R.E.CTRL.INST ( 20 ) /= V_E_CTRL_INST20_shadow_intermed_1) else '0';
dfp_trap_vector(156) <= '1' when (R.E.CTRL.INST ( 20 ) /= DE_INST20_shadow_intermed_3) else '0';
dfp_trap_vector(157) <= '1' when (R.E.CTRL.INST ( 20 ) /= V_A_CTRL_INST20_shadow_intermed_3) else '0';
dfp_trap_vector(158) <= '1' when (R.E.CTRL.INST ( 20 ) /= RIN_E_CTRL_INST20_intermed_2) else '0';
dfp_trap_vector(159) <= '1' when (R.E.CTRL.INST ( 20 ) /= R_A_CTRL_INST20_intermed_2) else '0';
dfp_trap_vector(160) <= '1' when (R.X.DATA ( 0 ) ( 0 ) /= RIN_X_DATA00_intermed_2) else '0';
dfp_trap_vector(161) <= '1' when (R.X.DATA ( 0 ) ( 0 ) /= V_X_DATA00_shadow_intermed_1) else '0';
dfp_trap_vector(162) <= '1' when (R.X.DATA ( 0 ) ( 0 ) /= DCO_DATA00_intermed_2) else '0';
dfp_trap_vector(163) <= '1' when (R.X.DATA ( 0 ) ( 0 ) /= V_X_DATA00_shadow_intermed_2) else '0';
dfp_trap_vector(164) <= '1' when (R.X.DATA ( 0 ) ( 0 ) /= RIN_X_DATA00_intermed_1) else '0';
dfp_trap_vector(165) <= '1' when (R.X.DATA ( 0 ) ( 0 ) /= V_X_DATA00_shadow_intermed_2) else '0';
dfp_trap_vector(166) <= '1' when (R.X.DATA ( 0 ) ( 0 ) /= R_X_DATA00_intermed_2) else '0';
dfp_trap_vector(167) <= '1' when (R.X.DATA ( 0 ) ( 0 ) /= RIN_X_DATA00_intermed_2) else '0';
dfp_trap_vector(168) <= '1' when (R.X.DATA ( 0 ) ( 0 ) /= R_X_DATA00_intermed_2) else '0';
dfp_trap_vector(169) <= '1' when (R.X.DATA ( 0 ) ( 4 DOWNTO 0 ) /= RIN_X_DATA04DOWNTO0_intermed_1) else '0';
dfp_trap_vector(170) <= '1' when (R.X.DATA ( 0 ) ( 4 DOWNTO 0 ) /= V_X_DATA04DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(171) <= '1' when (R.X.DATA ( 0 ) ( 4 DOWNTO 0 ) /= R_X_DATA04DOWNTO0_intermed_2) else '0';
dfp_trap_vector(172) <= '1' when (R.X.DATA ( 0 ) ( 4 DOWNTO 0 ) /= R_X_DATA04DOWNTO0_intermed_2) else '0';
dfp_trap_vector(173) <= '1' when (R.X.DATA ( 0 ) ( 4 DOWNTO 0 ) /= V_X_DATA04DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(174) <= '1' when (R.X.DATA ( 0 ) ( 4 DOWNTO 0 ) /= DCO_DATA04DOWNTO0_intermed_2) else '0';
dfp_trap_vector(175) <= '1' when (R.X.DATA ( 0 ) ( 4 DOWNTO 0 ) /= RIN_X_DATA04DOWNTO0_intermed_2) else '0';
dfp_trap_vector(176) <= '1' when (R.X.DATA ( 0 ) ( 4 DOWNTO 0 ) /= RIN_X_DATA04DOWNTO0_intermed_2) else '0';
dfp_trap_vector(177) <= '1' when (R.X.DATA ( 0 ) ( 4 DOWNTO 0 ) /= V_X_DATA04DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(178) <= '1' when (RFI.REN1 /= DCO.SCANEN) else '0';
dfp_trap_vector(179) <= '1' when (RFI.REN1 /= RIN_A_RFE1_intermed_1) else '0';
dfp_trap_vector(180) <= '1' when (RFI.REN1 /= DE_REN1_shadow) else '0';
dfp_trap_vector(181) <= '1' when (RFI.REN1 /= V_A_RFE1_shadow_intermed_1) else '0';
dfp_trap_vector(182) <= '1' when (RFI.REN1 /= R.A.RFE1) else '0';
dfp_trap_vector(183) <= '1' when (RFI.REN1 /= '1') else '0';
dfp_trap_vector(184) <= '1' when (RFI.REN2 /= DCO.SCANEN) else '0';
dfp_trap_vector(185) <= '1' when (RFI.REN2 /= RIN_A_RFE2_intermed_1) else '0';
dfp_trap_vector(186) <= '1' when (RFI.REN2 /= V_A_RFE2_shadow_intermed_1) else '0';
dfp_trap_vector(187) <= '1' when (RFI.REN2 /= DE_REN2_shadow) else '0';
dfp_trap_vector(188) <= '1' when (RFI.REN2 /= R.A.RFE2) else '0';
dfp_trap_vector(189) <= '1' when (RFI.DIAG(0) /= DCO.TESTEN) else '0';
dfp_trap_vector(190) <= '1' when (RFI.DIAG /= "0000") else '0';
dfp_trap_vector(191) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= R_M_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(192) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= RIN_M_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(193) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_6) else '0';
dfp_trap_vector(194) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= RIN_A_CTRL_PC31DOWNTO2_intermed_7) else '0';
dfp_trap_vector(195) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= R_A_CTRL_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(196) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(197) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= R_X_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(198) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= V_D_PC31DOWNTO2_shadow_intermed_8) else '0';
dfp_trap_vector(199) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(200) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= RIN_D_PC31DOWNTO2_intermed_8) else '0';
dfp_trap_vector(201) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_2) else '0';
dfp_trap_vector(202) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= V_F_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(203) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= V_F_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(204) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= RIN_F_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(205) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= RIN_X_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(206) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= IRIN_ADDR31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(207) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= R_E_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(208) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_7) else '0';
dfp_trap_vector(209) <= '1' when (R.F.PC ( 2 DOWNTO 2 ) /= "1") else '0';
dfp_trap_vector(210) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(211) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= R_D_PC31DOWNTO2_intermed_7) else '0';
dfp_trap_vector(212) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= RIN_F_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(213) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= IR_ADDR31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(214) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= RIN_E_CTRL_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(215) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= R_F_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(216) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= V_X_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(217) <= '1' when (R.F.PC ( 31 DOWNTO 2 ) /= VIR_ADDR31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(218) <= '1' when (ICI.DPC(31 downto 2) /= V_D_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(219) <= '1' when (ICI.DPC(31 downto 2) /= RIN_D_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(220) <= '1' when (ICI.DPC /= x"00000000") else '0';
dfp_trap_vector(221) <= '1' when (ICI.DPC(31 downto 2) /= R.D.PC ( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(222) <= '1' when (ICI.DPC(31 downto 2) /= R_D_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(223) <= '1' when (ICI.DPC(31 downto 2) /= V_D_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(224) <= '1' when (ICI.DPC(31 downto 2) /= RIN_D_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(225) <= '1' when (R.D.PC ( 31 DOWNTO 2 ) /= V_D_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(226) <= '1' when (R.D.PC ( 31 DOWNTO 2 ) /= RIN_D_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(227) <= '1' when (R.D.PC ( 31 DOWNTO 2 ) /= R_D_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(228) <= '1' when (R.D.PC ( 31 DOWNTO 2 ) /= V_D_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(229) <= '1' when (R.D.PC ( 31 DOWNTO 2 ) /= RIN_D_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(230) <= '1' when (ICI.FPC(31 downto 2) /= R_M_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(231) <= '1' when (ICI.FPC(31 downto 2) /= RIN_M_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(232) <= '1' when (ICI.FPC(31 downto 2) /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(233) <= '1' when (ICI.FPC(31 downto 2) /= RIN_A_CTRL_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(234) <= '1' when (ICI.FPC(31 downto 2) /= R_A_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(235) <= '1' when (ICI.FPC(31 downto 2) /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(236) <= '1' when (ICI.FPC(31 downto 2) /= R_X_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(237) <= '1' when (ICI.FPC(31 downto 2) /= V_D_PC31DOWNTO2_shadow_intermed_7) else '0';
dfp_trap_vector(238) <= '1' when (ICI.FPC(31 downto 2) /= XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(239) <= '1' when (ICI.FPC(31 downto 2) /= RIN_D_PC31DOWNTO2_intermed_7) else '0';
dfp_trap_vector(240) <= '1' when (ICI.FPC(31 downto 2) /= EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_2) else '0';
dfp_trap_vector(241) <= '1' when (ICI.FPC(31 downto 2) /= V_F_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(242) <= '1' when (ICI.FPC(31 downto 2) /= V_F_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(243) <= '1' when (ICI.FPC(31 downto 2) /= RIN_F_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(244) <= '1' when (ICI.FPC(31 downto 2) /= RIN_X_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(245) <= '1' when (ICI.FPC /= X"00000000") else '0';
dfp_trap_vector(246) <= '1' when (ICI.FPC(31 downto 2) /= IRIN_ADDR31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(247) <= '1' when (ICI.FPC(31 downto 2) /= R_E_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(248) <= '1' when (ICI.FPC(31 downto 2) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_6) else '0';
dfp_trap_vector(249) <= '1' when (ICI.FPC(0) /= '1') else '0';
dfp_trap_vector(250) <= '1' when (ICI.FPC(31 downto 2) /= EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(251) <= '1' when (ICI.FPC(31 downto 2) /= R_D_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(252) <= '1' when (ICI.FPC(31 downto 2) /= R.F.PC ( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(253) <= '1' when (ICI.FPC(31 downto 2) /= RIN_F_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(254) <= '1' when (ICI.FPC(31 downto 2) /= IR_ADDR31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(255) <= '1' when (ICI.FPC(31 downto 2) /= RIN_E_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(256) <= '1' when (ICI.FPC(31 downto 2) /= R_F_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(257) <= '1' when (ICI.FPC(31 downto 2) /= V_X_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(258) <= '1' when (ICI.FPC(31 downto 2) /= VIR_ADDR31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(259) <= '1' when (ICI.RPC(31 downto 2) /= R_M_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(260) <= '1' when (ICI.RPC(31 downto 2) /= RIN_M_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(261) <= '1' when (ICI.RPC(31 downto 2) /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(262) <= '1' when (ICI.RPC(31 downto 2) /= RIN_A_CTRL_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(263) <= '1' when (ICI.RPC(31 downto 2) /= R_A_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(264) <= '1' when (ICI.RPC(31 downto 2) /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(265) <= '1' when (ICI.RPC(31 downto 2) /= NPC31DOWNTO2_shadow) else '0';
dfp_trap_vector(266) <= '1' when (ICI.RPC(31 downto 2) /= R_X_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(267) <= '1' when (ICI.RPC(31 downto 2) /= V_D_PC31DOWNTO2_shadow_intermed_7) else '0';
dfp_trap_vector(268) <= '1' when (ICI.RPC(31 downto 2) /= XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(269) <= '1' when (ICI.RPC(31 downto 2) /= RIN_D_PC31DOWNTO2_intermed_7) else '0';
dfp_trap_vector(270) <= '1' when (ICI.RPC(31 downto 2) /= EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_1) else '0';
dfp_trap_vector(271) <= '1' when (ICI.RPC(31 downto 2) /= V_F_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(272) <= '1' when (ICI.RPC(31 downto 2) /= RIN_F_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(273) <= '1' when (ICI.RPC(31 downto 2) /= RIN_X_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(274) <= '1' when (ICI.RPC /= X"00000000") else '0';
dfp_trap_vector(275) <= '1' when (ICI.RPC(31 downto 2) /= IRIN_ADDR31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(276) <= '1' when (ICI.RPC(31 downto 2) /= R_E_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(277) <= '1' when (ICI.RPC(31 downto 2) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_6) else '0';
dfp_trap_vector(278) <= '1' when (ICI.RPC(31 downto 2) /= EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(279) <= '1' when (ICI.RPC(31 downto 2) /= R_D_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(280) <= '1' when (ICI.RPC(31 downto 2) /= IR_ADDR31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(281) <= '1' when (ICI.RPC(31 downto 2) /= RIN_E_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(282) <= '1' when (ICI.RPC(31 downto 2) /= R.F.PC( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(283) <= '1' when (ICI.RPC(31 downto 2) /= V_X_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(284) <= '1' when (ICI.RPC(31 downto 2) /= VIR_ADDR31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(285) <= '1' when (ICI.FLUSHL /= '0') else '0';
dfp_trap_vector(286) <= '1' when (MULI.START /= R.A.MULSTART) else '0';
dfp_trap_vector(287) <= '1' when (MULI.START /= V_X_ANNUL_ALL_shadow_intermed_1) else '0';
dfp_trap_vector(288) <= '1' when (MULI.START /= RIN_A_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(289) <= '1' when (MULI.START /= R.A.CTRL.ANNUL) else '0';
dfp_trap_vector(290) <= '1' when (MULI.START /= V_A_MULSTART_shadow_intermed_1) else '0';
dfp_trap_vector(291) <= '1' when (MULI.START /= RIN_X_ANNUL_ALL_intermed_2) else '0';
dfp_trap_vector(292) <= '1' when (MULI.START /= R_X_ANNUL_ALL_intermed_1) else '0';
dfp_trap_vector(293) <= '1' when (MULI.START /= RIN_A_MULSTART_intermed_1) else '0';
dfp_trap_vector(294) <= '1' when (MULI.START /= '1') else '0';
dfp_trap_vector(295) <= '1' when (MULI.START /= '0') else '0';
dfp_trap_vector(296) <= '1' when (MULI.START /= V_A_CTRL_ANNUL_shadow_intermed_1) else '0';
dfp_trap_vector(297) <= '1' when (MULI.OP1(31) /= RIN_X_DATA031_intermed_1) else '0';
dfp_trap_vector(298) <= '1' when (MULI.OP1(31 downto 0) /= V_X_DATA0_shadow_intermed_2) else '0';
dfp_trap_vector(299) <= '1' when (MULI.OP1(19) /= DE_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(300) <= '1' when (MULI.OP1(31) /= RIN_E_OP131_intermed_1) else '0';
dfp_trap_vector(301) <= '1' when (MULI.OP1(19) /= V_A_CTRL_INST19_shadow_intermed_3) else '0';
dfp_trap_vector(302) <= '1' when (MULI.OP1(31 downto 0) /= RIN_X_DATA0_intermed_1) else '0';
dfp_trap_vector(303) <= '1' when (MULI.OP1(31) /= V_E_OP131_shadow_intermed_1) else '0';
dfp_trap_vector(304) <= '1' when (MULI.OP1(31) /= V_X_DATA031_shadow_intermed_1) else '0';
dfp_trap_vector(305) <= '1' when (MULI.OP1(31) /= R.E.OP1( 31 )) else '0';
dfp_trap_vector(306) <= '1' when (MULI.OP1(19) /= V_E_CTRL_INST19_shadow_intermed_1) else '0';
dfp_trap_vector(307) <= '1' when (MULI.OP1(31 downto 0) /= V_E_OP1_shadow_intermed_1) else '0';
dfp_trap_vector(308) <= '1' when (MULI.OP1(31) /= V_X_DATA031_shadow_intermed_2) else '0';
dfp_trap_vector(309) <= '1' when (MULI.OP1(19) /= V_E_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(310) <= '1' when (MULI.OP1(31) /= RIN_X_DATA031_intermed_2) else '0';
dfp_trap_vector(311) <= '1' when (MULI.OP1(31 downto 0) /= RIN_E_OP1_intermed_1) else '0';
dfp_trap_vector(312) <= '1' when (MULI.OP1(19) /= R_E_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(313) <= '1' when (MULI.OP1(31 downto 0) /= V_X_DATA0_shadow_intermed_1) else '0';
dfp_trap_vector(314) <= '1' when (MULI.OP1(31 downto 0) /= EX_OP1_shadow) else '0';
dfp_trap_vector(315) <= '1' when (MULI.OP1(31) /= DCO_DATA031_intermed_1) else '0';
dfp_trap_vector(316) <= '1' when (MULI.OP1(31) /= R_X_DATA031_intermed_1) else '0';
dfp_trap_vector(317) <= '1' when (MULI.OP1(31) /= EX_OP131_shadow) else '0';
dfp_trap_vector(318) <= '1' when (MULI.OP1(19) /= RIN_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(319) <= '1' when (MULI.OP1(31 downto 0) /= R_X_DATA0_intermed_1) else '0';
dfp_trap_vector(320) <= '1' when (MULI.OP1(31 downto 0) /= R.X.DATA ( 0 )) else '0';
dfp_trap_vector(321) <= '1' when (MULI.OP1(19) /= R_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(322) <= '1' when (MULI.OP1(19) /= R_A_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(323) <= '1' when (MULI.OP1(19) /= RIN_A_CTRL_INST19_intermed_3) else '0';
dfp_trap_vector(324) <= '1' when (MULI.OP1(19) /= RIN_E_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(325) <= '1' when (MULI.OP1(19) /= R.E.CTRL.INST ( 19 )) else '0';
dfp_trap_vector(326) <= '1' when (MULI.OP1(31) /= R.X.DATA ( 0 )( 31 )) else '0';
dfp_trap_vector(327) <= '1' when (MULI.OP1(31 downto 0) /= DCO_DATA0_intermed_1) else '0';
dfp_trap_vector(328) <= '1' when (MULI.OP1(31 downto 0) /= RIN_X_DATA0_intermed_2) else '0';
dfp_trap_vector(329) <= '1' when (MULI.OP1(19) /= RIN_E_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(330) <= '1' when (MULI.OP1(31 downto 0) /= R.E.OP1) else '0';
dfp_trap_vector(331) <= '1' when (MULI.OP1(19) /= V_A_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(332) <= '1' when (MULI.OP2(31) /= RIN_X_DATA031_intermed_1) else '0';
dfp_trap_vector(333) <= '1' when (MULI.OP2(31 downto 0) /= V_X_DATA0_shadow_intermed_2) else '0';
dfp_trap_vector(334) <= '1' when (MULI.OP2(19) /= DE_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(335) <= '1' when (MULI.OP2(31 downto 0) /= MUL_OP2_shadow) else '0';
dfp_trap_vector(336) <= '1' when (MULI.OP2(19) /= V_A_CTRL_INST19_shadow_intermed_3) else '0';
dfp_trap_vector(337) <= '1' when (MULI.OP2(31 downto 0) /= RIN_X_DATA0_intermed_1) else '0';
dfp_trap_vector(338) <= '1' when (MULI.OP2(31) /= V_X_DATA031_shadow_intermed_1) else '0';
dfp_trap_vector(339) <= '1' when (MULI.OP2(19) /= V_E_CTRL_INST19_shadow_intermed_1) else '0';
dfp_trap_vector(340) <= '1' when (MULI.OP2(31) /= V_X_DATA031_shadow_intermed_2) else '0';
dfp_trap_vector(341) <= '1' when (MULI.OP2(31 downto 0) /= V_E_OP2_shadow_intermed_1) else '0';
dfp_trap_vector(342) <= '1' when (MULI.OP2(31 downto 0) /= RIN_E_OP2_intermed_1) else '0';
dfp_trap_vector(343) <= '1' when (MULI.OP2(19) /= V_E_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(344) <= '1' when (MULI.OP2(31) /= RIN_X_DATA031_intermed_2) else '0';
dfp_trap_vector(345) <= '1' when (MULI.OP2(31) /= EX_OP231_shadow) else '0';
dfp_trap_vector(346) <= '1' when (MULI.OP2(19) /= R_E_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(347) <= '1' when (MULI.OP2(31 downto 0) /= V_X_DATA0_shadow_intermed_1) else '0';
dfp_trap_vector(348) <= '1' when (MULI.OP2(31 downto 0) /= EX_OP2_shadow) else '0';
dfp_trap_vector(349) <= '1' when (MULI.OP2(31) /= DCO_DATA031_intermed_1) else '0';
dfp_trap_vector(350) <= '1' when (MULI.OP2(31) /= R_X_DATA031_intermed_1) else '0';
dfp_trap_vector(351) <= '1' when (MULI.OP2(19) /= RIN_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(352) <= '1' when (MULI.OP2(31 downto 0) /= R_X_DATA0_intermed_1) else '0';
dfp_trap_vector(353) <= '1' when (MULI.OP2(31 downto 0) /= R.X.DATA ( 0 )) else '0';
dfp_trap_vector(354) <= '1' when (MULI.OP2(19) /= R_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(355) <= '1' when (MULI.OP2(31) /= RIN_E_OP231_intermed_1) else '0';
dfp_trap_vector(356) <= '1' when (MULI.OP2(31) /= R.E.OP2( 31 )) else '0';
dfp_trap_vector(357) <= '1' when (MULI.OP2(31) /= MUL_OP231_shadow) else '0';
dfp_trap_vector(358) <= '1' when (MULI.OP2(19) /= R_A_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(359) <= '1' when (MULI.OP2(19) /= RIN_A_CTRL_INST19_intermed_3) else '0';
dfp_trap_vector(360) <= '1' when (MULI.OP2(19) /= RIN_E_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(361) <= '1' when (MULI.OP2(31 downto 0) /= R.E.OP2) else '0';
dfp_trap_vector(362) <= '1' when (MULI.OP2(19) /= R.E.CTRL.INST ( 19 )) else '0';
dfp_trap_vector(363) <= '1' when (MULI.OP2(31) /= V_E_OP231_shadow_intermed_1) else '0';
dfp_trap_vector(364) <= '1' when (MULI.OP2(31) /= R.X.DATA ( 0 )( 31 )) else '0';
dfp_trap_vector(365) <= '1' when (MULI.OP2(31 downto 0) /= DCO_DATA0_intermed_1) else '0';
dfp_trap_vector(366) <= '1' when (MULI.OP2(31 downto 0) /= RIN_X_DATA0_intermed_2) else '0';
dfp_trap_vector(367) <= '1' when (MULI.OP2(19) /= RIN_E_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(368) <= '1' when (MULI.OP2(19) /= V_A_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(369) <= '1' when (R.E.CTRL.INST ( 24 ) /= V_A_CTRL_INST24_shadow_intermed_3) else '0';
dfp_trap_vector(370) <= '1' when (R.E.CTRL.INST ( 24 ) /= V_E_CTRL_INST24_shadow_intermed_2) else '0';
dfp_trap_vector(371) <= '1' when (R.E.CTRL.INST ( 24 ) /= DE_INST24_shadow_intermed_3) else '0';
dfp_trap_vector(372) <= '1' when (R.E.CTRL.INST ( 24 ) /= V_E_CTRL_INST24_shadow_intermed_1) else '0';
dfp_trap_vector(373) <= '1' when (R.E.CTRL.INST ( 24 ) /= R_A_CTRL_INST24_intermed_2) else '0';
dfp_trap_vector(374) <= '1' when (R.E.CTRL.INST ( 24 ) /= RIN_A_CTRL_INST24_intermed_2) else '0';
dfp_trap_vector(375) <= '1' when (R.E.CTRL.INST ( 24 ) /= V_A_CTRL_INST24_shadow_intermed_2) else '0';
dfp_trap_vector(376) <= '1' when (R.E.CTRL.INST ( 24 ) /= RIN_A_CTRL_INST24_intermed_3) else '0';
dfp_trap_vector(377) <= '1' when (R.E.CTRL.INST ( 24 ) /= RIN_E_CTRL_INST24_intermed_2) else '0';
dfp_trap_vector(378) <= '1' when (R.E.CTRL.INST ( 24 ) /= R_E_CTRL_INST24_intermed_2) else '0';
dfp_trap_vector(379) <= '1' when (R.E.CTRL.INST ( 24 ) /= R_A_CTRL_INST24_intermed_1) else '0';
dfp_trap_vector(380) <= '1' when (R.E.CTRL.INST ( 24 ) /= RIN_E_CTRL_INST24_intermed_1) else '0';
dfp_trap_vector(381) <= '1' when (DIVI.START /= R.A.DIVSTART) else '0';
dfp_trap_vector(382) <= '1' when (DIVI.START /= V_X_ANNUL_ALL_shadow_intermed_1) else '0';
dfp_trap_vector(383) <= '1' when (DIVI.START /= RIN_A_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(384) <= '1' when (DIVI.START /= R.A.CTRL.ANNUL) else '0';
dfp_trap_vector(385) <= '1' when (DIVI.START /= RIN_A_DIVSTART_intermed_1) else '0';
dfp_trap_vector(386) <= '1' when (DIVI.START /= RIN_X_ANNUL_ALL_intermed_2) else '0';
dfp_trap_vector(387) <= '1' when (DIVI.START /= R_X_ANNUL_ALL_intermed_1) else '0';
dfp_trap_vector(388) <= '1' when (DIVI.START /= V_A_DIVSTART_shadow_intermed_1) else '0';
dfp_trap_vector(389) <= '1' when (DIVI.START /= '1') else '0';
dfp_trap_vector(390) <= '1' when (DIVI.START /= '0') else '0';
dfp_trap_vector(391) <= '1' when (DIVI.START /= V_A_CTRL_ANNUL_shadow_intermed_1) else '0';
dfp_trap_vector(392) <= '1' when (DIVI.OP1(31) /= RIN_X_DATA031_intermed_1) else '0';
dfp_trap_vector(393) <= '1' when (DIVI.OP1(31 downto 0) /= V_X_DATA0_shadow_intermed_2) else '0';
dfp_trap_vector(394) <= '1' when (DIVI.OP1(19) /= DE_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(395) <= '1' when (DIVI.OP1(31) /= RIN_E_OP131_intermed_1) else '0';
dfp_trap_vector(396) <= '1' when (DIVI.OP1(19) /= V_A_CTRL_INST19_shadow_intermed_3) else '0';
dfp_trap_vector(397) <= '1' when (DIVI.OP1(31 downto 0) /= RIN_X_DATA0_intermed_1) else '0';
dfp_trap_vector(398) <= '1' when (DIVI.OP1(31) /= V_E_OP131_shadow_intermed_1) else '0';
dfp_trap_vector(399) <= '1' when (DIVI.OP1(31) /= V_X_DATA031_shadow_intermed_1) else '0';
dfp_trap_vector(400) <= '1' when (DIVI.OP1(31) /= R.E.OP1( 31 )) else '0';
dfp_trap_vector(401) <= '1' when (DIVI.OP1(19) /= V_E_CTRL_INST19_shadow_intermed_1) else '0';
dfp_trap_vector(402) <= '1' when (DIVI.OP1(31 downto 0) /= V_E_OP1_shadow_intermed_1) else '0';
dfp_trap_vector(403) <= '1' when (DIVI.OP1(31) /= V_X_DATA031_shadow_intermed_2) else '0';
dfp_trap_vector(404) <= '1' when (DIVI.OP1(19) /= V_E_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(405) <= '1' when (DIVI.OP1(31) /= RIN_X_DATA031_intermed_2) else '0';
dfp_trap_vector(406) <= '1' when (DIVI.OP1(31 downto 0) /= RIN_E_OP1_intermed_1) else '0';
dfp_trap_vector(407) <= '1' when (DIVI.OP1(19) /= R_E_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(408) <= '1' when (DIVI.OP1(31 downto 0) /= V_X_DATA0_shadow_intermed_1) else '0';
dfp_trap_vector(409) <= '1' when (DIVI.OP1(31 downto 0) /= EX_OP1_shadow) else '0';
dfp_trap_vector(410) <= '1' when (DIVI.OP1(31) /= DCO_DATA031_intermed_1) else '0';
dfp_trap_vector(411) <= '1' when (DIVI.OP1(31) /= R_X_DATA031_intermed_1) else '0';
dfp_trap_vector(412) <= '1' when (DIVI.OP1(31) /= EX_OP131_shadow) else '0';
dfp_trap_vector(413) <= '1' when (DIVI.OP1(19) /= RIN_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(414) <= '1' when (DIVI.OP1(31 downto 0) /= R_X_DATA0_intermed_1) else '0';
dfp_trap_vector(415) <= '1' when (DIVI.OP1(31 downto 0) /= R.X.DATA ( 0 )) else '0';
dfp_trap_vector(416) <= '1' when (DIVI.OP1(19) /= R_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(417) <= '1' when (DIVI.OP1(19) /= R_A_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(418) <= '1' when (DIVI.OP1(19) /= RIN_A_CTRL_INST19_intermed_3) else '0';
dfp_trap_vector(419) <= '1' when (DIVI.OP1(19) /= RIN_E_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(420) <= '1' when (DIVI.OP1(19) /= R.E.CTRL.INST ( 19 )) else '0';
dfp_trap_vector(421) <= '1' when (DIVI.OP1(31) /= R.X.DATA ( 0 )( 31 )) else '0';
dfp_trap_vector(422) <= '1' when (DIVI.OP1(31 downto 0) /= DCO_DATA0_intermed_1) else '0';
dfp_trap_vector(423) <= '1' when (DIVI.OP1(31 downto 0) /= RIN_X_DATA0_intermed_2) else '0';
dfp_trap_vector(424) <= '1' when (DIVI.OP1(19) /= RIN_E_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(425) <= '1' when (DIVI.OP1(31 downto 0) /= R.E.OP1) else '0';
dfp_trap_vector(426) <= '1' when (DIVI.OP1(19) /= V_A_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(427) <= '1' when (DIVI.OP2(31) /= RIN_X_DATA031_intermed_1) else '0';
dfp_trap_vector(428) <= '1' when (DIVI.OP2(31 downto 0) /= V_X_DATA0_shadow_intermed_2) else '0';
dfp_trap_vector(429) <= '1' when (DIVI.OP2(19) /= DE_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(430) <= '1' when (DIVI.OP2(19) /= V_A_CTRL_INST19_shadow_intermed_3) else '0';
dfp_trap_vector(431) <= '1' when (DIVI.OP2(31 downto 0) /= RIN_X_DATA0_intermed_1) else '0';
dfp_trap_vector(432) <= '1' when (DIVI.OP2(31) /= V_X_DATA031_shadow_intermed_1) else '0';
dfp_trap_vector(433) <= '1' when (DIVI.OP2(31) /= EX_OP231_shadow) else '0';
dfp_trap_vector(434) <= '1' when (DIVI.OP2(19) /= V_E_CTRL_INST19_shadow_intermed_1) else '0';
dfp_trap_vector(435) <= '1' when (DIVI.OP2(31) /= V_X_DATA031_shadow_intermed_2) else '0';
dfp_trap_vector(436) <= '1' when (DIVI.OP2(31 downto 0) /= V_E_OP2_shadow_intermed_1) else '0';
dfp_trap_vector(437) <= '1' when (DIVI.OP2(31 downto 0) /= RIN_E_OP2_intermed_1) else '0';
dfp_trap_vector(438) <= '1' when (DIVI.OP2(19) /= V_E_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(439) <= '1' when (DIVI.OP2(31) /= RIN_X_DATA031_intermed_2) else '0';
dfp_trap_vector(440) <= '1' when (DIVI.OP2(19) /= R_E_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(441) <= '1' when (DIVI.OP2(31 downto 0) /= V_X_DATA0_shadow_intermed_1) else '0';
dfp_trap_vector(442) <= '1' when (DIVI.OP2(31 downto 0) /= EX_OP2_shadow) else '0';
dfp_trap_vector(443) <= '1' when (DIVI.OP2(31) /= DCO_DATA031_intermed_1) else '0';
dfp_trap_vector(444) <= '1' when (DIVI.OP2(31) /= R_X_DATA031_intermed_1) else '0';
dfp_trap_vector(445) <= '1' when (DIVI.OP2(19) /= RIN_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(446) <= '1' when (DIVI.OP2(31 downto 0) /= R_X_DATA0_intermed_1) else '0';
dfp_trap_vector(447) <= '1' when (DIVI.OP2(31 downto 0) /= R.X.DATA ( 0 )) else '0';
dfp_trap_vector(448) <= '1' when (DIVI.OP2(19) /= R_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(449) <= '1' when (DIVI.OP2(31) /= RIN_E_OP231_intermed_1) else '0';
dfp_trap_vector(450) <= '1' when (DIVI.OP2(31) /= R.E.OP2( 31 )) else '0';
dfp_trap_vector(451) <= '1' when (DIVI.OP2(19) /= R_A_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(452) <= '1' when (DIVI.OP2(19) /= RIN_A_CTRL_INST19_intermed_3) else '0';
dfp_trap_vector(453) <= '1' when (DIVI.OP2(19) /= RIN_E_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(454) <= '1' when (DIVI.OP2(31 downto 0) /= R.E.OP2) else '0';
dfp_trap_vector(455) <= '1' when (DIVI.OP2(19) /= R.E.CTRL.INST ( 19 )) else '0';
dfp_trap_vector(456) <= '1' when (DIVI.OP2(31) /= V_E_OP231_shadow_intermed_1) else '0';
dfp_trap_vector(457) <= '1' when (DIVI.OP2(31) /= R.X.DATA ( 0 )( 31 )) else '0';
dfp_trap_vector(458) <= '1' when (DIVI.OP2(31 downto 0) /= DCO_DATA0_intermed_1) else '0';
dfp_trap_vector(459) <= '1' when (DIVI.OP2(31 downto 0) /= RIN_X_DATA0_intermed_2) else '0';
dfp_trap_vector(460) <= '1' when (DIVI.OP2(19) /= RIN_E_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(461) <= '1' when (DIVI.OP2(19) /= V_A_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(462) <= '1' when (R.A.CTRL.INST ( 19 ) /= DE_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(463) <= '1' when (R.A.CTRL.INST ( 19 ) /= V_A_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(464) <= '1' when (R.A.CTRL.INST ( 19 ) /= RIN_A_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(465) <= '1' when (R.A.CTRL.INST ( 19 ) /= R_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(466) <= '1' when (R.A.CTRL.INST ( 19 ) /= RIN_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(467) <= '1' when (R.A.CTRL.INST ( 19 ) /= V_A_CTRL_INST19_shadow_intermed_1) else '0';
dfp_trap_vector(468) <= '1' when (DIVI.Y(19) /= DE_INST19_shadow_intermed_1) else '0';
dfp_trap_vector(469) <= '1' when (DIVI.Y(31) /= RIN_M_Y31_intermed_1) else '0';
dfp_trap_vector(470) <= '1' when (DIVI.Y(31 downto 0) /= RIN_M_Y_intermed_1) else '0';
dfp_trap_vector(471) <= '1' when (DIVI.Y(19) /= V_A_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(472) <= '1' when (DIVI.Y(19) /= V_E_CTRL_INST19_shadow_intermed_1) else '0';
dfp_trap_vector(473) <= '1' when (DIVI.Y(31) /= V_M_Y31_shadow_intermed_2) else '0';
dfp_trap_vector(474) <= '1' when (DIVI.Y(31 downto 0) /= V_M_Y_shadow_intermed_1) else '0';
dfp_trap_vector(475) <= '1' when (DIVI.Y(19) /= V_E_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(476) <= '1' when (DIVI.Y(31 downto 0) /= R.M.Y) else '0';
dfp_trap_vector(477) <= '1' when (DIVI.Y(19) /= R_E_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(478) <= '1' when (DIVI.Y(31) /= V_M_Y31_shadow_intermed_1) else '0';
dfp_trap_vector(479) <= '1' when (DIVI.Y(19) /= RIN_A_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(480) <= '1' when (DIVI.Y(0) /= DSIGN_shadow) else '0';
dfp_trap_vector(481) <= '1' when (DIVI.Y(31) /= RIN_M_Y31_intermed_2) else '0';
dfp_trap_vector(482) <= '1' when (DIVI.Y(19) /= R_A_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(483) <= '1' when (DIVI.Y(31) /= R_M_Y31_intermed_1) else '0';
dfp_trap_vector(484) <= '1' when (DIVI.Y(19) /= R.A.CTRL.INST ( 19 )) else '0';
dfp_trap_vector(485) <= '1' when (DIVI.Y(19) /= RIN_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(486) <= '1' when (DIVI.Y(19) /= RIN_E_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(487) <= '1' when (DIVI.Y(19) /= R.E.CTRL.INST ( 19 )) else '0';
dfp_trap_vector(488) <= '1' when (DIVI.Y(31) /= R.M.Y ( 31 )) else '0';
dfp_trap_vector(489) <= '1' when (DIVI.Y(19) /= RIN_E_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(490) <= '1' when (DIVI.Y(19) /= V_A_CTRL_INST19_shadow_intermed_1) else '0';
dfp_trap_vector(491) <= '1' when (R.M.Y ( 31 ) /= RIN_M_Y31_intermed_1) else '0';
dfp_trap_vector(492) <= '1' when (R.M.Y ( 31 ) /= V_M_Y31_shadow_intermed_2) else '0';
dfp_trap_vector(493) <= '1' when (R.M.Y ( 31 ) /= V_M_Y31_shadow_intermed_1) else '0';
dfp_trap_vector(494) <= '1' when (R.M.Y ( 31 ) /= RIN_M_Y31_intermed_2) else '0';
dfp_trap_vector(495) <= '1' when (R.M.Y ( 31 ) /= R_M_Y31_intermed_2) else '0';
dfp_trap_vector(496) <= '1' when (DSUR.CRDY ( 2 ) /= VDSU_CRDY2_shadow_intermed_2) else '0';
dfp_trap_vector(497) <= '1' when (DSUR.CRDY ( 2 ) /= DSUIN_CRDY2_intermed_1) else '0';
dfp_trap_vector(498) <= '1' when (DSUR.CRDY ( 2 ) /= VDSU_CRDY2_shadow_intermed_1) else '0';
dfp_trap_vector(499) <= '1' when (DSUR.CRDY ( 2 ) /= DSUIN_CRDY2_intermed_2) else '0';
dfp_trap_vector(500) <= '1' when (DSUR.CRDY ( 2 ) /= DSUR_CRDY2_intermed_2) else '0';
dfp_trap_vector(501) <= '1' when (DBGO.ERROR /= VP_ERROR_shadow_intermed_2) else '0';
dfp_trap_vector(502) <= '1' when (DBGO.ERROR /= R.X.NERROR) else '0';
dfp_trap_vector(503) <= '1' when (DBGO.ERROR /= DUMMY) else '0';
dfp_trap_vector(504) <= '1' when (DBGO.ERROR /= RIN_X_NERROR_intermed_1) else '0';
dfp_trap_vector(505) <= '1' when (DBGO.ERROR /= '1') else '0';
dfp_trap_vector(506) <= '1' when (DBGO.ERROR /= '0') else '0';
dfp_trap_vector(507) <= '1' when (DBGO.ERROR /= RPIN_ERROR_intermed_2) else '0';
dfp_trap_vector(508) <= '1' when (DBGO.ERROR /= V_X_NERROR_shadow_intermed_1) else '0';
dfp_trap_vector(509) <= '1' when (DBGO.ERROR /= RP_ERROR_intermed_1) else '0';
dfp_trap_vector(510) <= '1' when (R.A.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_A_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(511) <= '1' when (R.A.CTRL.PC ( 31 DOWNTO 2 ) /= R_A_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(512) <= '1' when (R.A.CTRL.PC ( 31 DOWNTO 2 ) /= V_D_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(513) <= '1' when (R.A.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_D_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(514) <= '1' when (R.A.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_A_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(515) <= '1' when (R.A.CTRL.PC ( 31 DOWNTO 2 ) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(516) <= '1' when (R.A.CTRL.PC ( 31 DOWNTO 2 ) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(517) <= '1' when (R.A.CTRL.PC ( 31 DOWNTO 2 ) /= R_D_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(518) <= '1' when (R.E.CTRL.PC ( 31 DOWNTO 2 ) /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(519) <= '1' when (R.E.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_A_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(520) <= '1' when (R.E.CTRL.PC ( 31 DOWNTO 2 ) /= R_A_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(521) <= '1' when (R.E.CTRL.PC ( 31 DOWNTO 2 ) /= R_A_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(522) <= '1' when (R.E.CTRL.PC ( 31 DOWNTO 2 ) /= V_D_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(523) <= '1' when (R.E.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_D_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(524) <= '1' when (R.E.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_E_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(525) <= '1' when (R.E.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_A_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(526) <= '1' when (R.E.CTRL.PC ( 31 DOWNTO 2 ) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(527) <= '1' when (R.E.CTRL.PC ( 31 DOWNTO 2 ) /= R_E_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(528) <= '1' when (R.E.CTRL.PC ( 31 DOWNTO 2 ) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(529) <= '1' when (R.E.CTRL.PC ( 31 DOWNTO 2 ) /= R_D_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(530) <= '1' when (R.E.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_E_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(531) <= '1' when (R.E.CTRL.PC ( 31 DOWNTO 2 ) /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(532) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= R_M_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(533) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_M_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(534) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(535) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_A_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(536) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(537) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= R_A_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(538) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(539) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= R_A_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(540) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= R_E_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(541) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= V_D_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(542) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_D_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(543) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_E_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(544) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_A_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(545) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_M_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(546) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(547) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= R_E_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(548) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(549) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= R_D_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(550) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_E_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(551) <= '1' when (R.M.CTRL.PC ( 31 DOWNTO 2 ) /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(552) <= '1' when (RIN.X.RESULT ( 6 DOWNTO 0 ) /= V_X_RESULT6DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(553) <= '1' when (RIN.X.RESULT ( 6 DOWNTO 0 ) /= RIN_X_RESULT6DOWNTO0_intermed_2) else '0';
dfp_trap_vector(554) <= '1' when (RIN.X.RESULT ( 6 DOWNTO 0 ) /= R_X_RESULT6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(555) <= '1' when (RIN.X.RESULT ( 6 DOWNTO 0 ) /= V_X_RESULT6DOWNTO0_shadow) else '0';
dfp_trap_vector(556) <= '1' when (RIN.X.RESULT ( 6 DOWNTO 0 ) /= R.X.RESULT ( 6 DOWNTO 0 )) else '0';
dfp_trap_vector(557) <= '1' when (RIN.X.DATA ( 0 ) /= V_X_DATA0_shadow_intermed_1) else '0';
dfp_trap_vector(558) <= '1' when (RIN.X.DATA ( 0 ) /= V_X_DATA0_shadow) else '0';
dfp_trap_vector(559) <= '1' when (RIN.X.DATA ( 0 ) /= R_X_DATA0_intermed_1) else '0';
dfp_trap_vector(560) <= '1' when (RIN.X.DATA ( 0 ) /= R.X.DATA ( 0 )) else '0';
dfp_trap_vector(561) <= '1' when (RIN.X.DATA ( 0 ) /= DCO.DATA ( 0 )) else '0';
dfp_trap_vector(562) <= '1' when (RIN.X.DATA ( 0 ) /= RIN_X_DATA0_intermed_2) else '0';
dfp_trap_vector(563) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= R_M_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(564) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_M_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(565) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(566) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_A_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(567) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(568) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= V_X_CTRL_PC31DOWNTO2_shadow) else '0';
dfp_trap_vector(569) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= R_A_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(570) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(571) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= R_A_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(572) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= R_E_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(573) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= R_X_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(574) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= V_D_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(575) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_D_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(576) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_E_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(577) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_A_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(578) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_M_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(579) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_X_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(580) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(581) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= R.X.CTRL.PC ( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(582) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= R_E_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(583) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(584) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= R_D_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(585) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= R.M.CTRL.PC ( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(586) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_E_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(587) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(588) <= '1' when (RIN.X.CTRL.PC ( 31 DOWNTO 2 ) /= V_X_CTRL_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(589) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= V_X_CTRL_TT3DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(590) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= R_M_CTRL_TT3DOWNTO0_intermed_2) else '0';
dfp_trap_vector(591) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= V_M_CTRL_TT3DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(592) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(593) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= R_X_RESULT6DOWNTO03DOWNTO0_intermed_2) else '0';
dfp_trap_vector(594) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= R_A_CTRL_TT3DOWNTO0_intermed_4) else '0';
dfp_trap_vector(595) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= RIN_A_CTRL_TT3DOWNTO0_intermed_5) else '0';
dfp_trap_vector(596) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_3) else '0';
dfp_trap_vector(597) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= V_A_CTRL_TT3DOWNTO0_shadow_intermed_5) else '0';
dfp_trap_vector(598) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2) else '0';
dfp_trap_vector(599) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= R_W_S_TT3DOWNTO0_intermed_1) else '0';
dfp_trap_vector(600) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= R_X_RESULT6DOWNTO03DOWNTO0_intermed_1) else '0';
dfp_trap_vector(601) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= R_E_CTRL_TT3DOWNTO0_intermed_3) else '0';
dfp_trap_vector(602) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(603) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= RIN_W_S_TT3DOWNTO0_intermed_2) else '0';
dfp_trap_vector(604) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= V_E_CTRL_TT3DOWNTO0_shadow_intermed_4) else '0';
dfp_trap_vector(605) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= RIN_M_CTRL_TT3DOWNTO0_intermed_3) else '0';
dfp_trap_vector(606) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= RIN_X_CTRL_TT3DOWNTO0_intermed_2) else '0';
dfp_trap_vector(607) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= V_W_S_TT3DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(608) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= R_X_CTRL_TT3DOWNTO0_intermed_1) else '0';
dfp_trap_vector(609) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= RIN_E_CTRL_TT3DOWNTO0_intermed_4) else '0';
dfp_trap_vector(610) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= R.W.S.TT ( 3 DOWNTO 0 )) else '0';
dfp_trap_vector(611) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= V_W_S_TT3DOWNTO0_shadow) else '0';
dfp_trap_vector(612) <= '1' when (RIN.W.S.TT ( 3 DOWNTO 0 ) /= XC_VECTT3DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(613) <= '1' when (RIN.M.RESULT ( 1 DOWNTO 0 ) /= V_M_RESULT1DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(614) <= '1' when (RIN.M.RESULT ( 1 DOWNTO 0 ) /= R.M.RESULT ( 1 DOWNTO 0 )) else '0';
dfp_trap_vector(615) <= '1' when (RIN.M.RESULT ( 1 DOWNTO 0 ) /= RIN_M_RESULT1DOWNTO0_intermed_2) else '0';
dfp_trap_vector(616) <= '1' when (RIN.M.RESULT ( 1 DOWNTO 0 ) /= V_M_RESULT1DOWNTO0_shadow) else '0';
dfp_trap_vector(617) <= '1' when (RIN.M.RESULT ( 1 DOWNTO 0 ) /= R_M_RESULT1DOWNTO0_intermed_1) else '0';
dfp_trap_vector(618) <= '1' when (RIN.X.DATA ( 0 ) ( 31 ) /= RIN_X_DATA031_intermed_2) else '0';
dfp_trap_vector(619) <= '1' when (RIN.X.DATA ( 0 ) ( 31 ) /= V_X_DATA031_shadow_intermed_1) else '0';
dfp_trap_vector(620) <= '1' when (RIN.X.DATA ( 0 ) ( 31 ) /= V_X_DATA031_shadow_intermed_1) else '0';
dfp_trap_vector(621) <= '1' when (RIN.X.DATA ( 0 ) ( 31 ) /= R.X.DATA ( 0 ) ( 31 )) else '0';
dfp_trap_vector(622) <= '1' when (RIN.X.DATA ( 0 ) ( 31 ) /= RIN_X_DATA031_intermed_2) else '0';
dfp_trap_vector(623) <= '1' when (RIN.X.DATA ( 0 ) ( 31 ) /= DCO_DATA031_intermed_1) else '0';
dfp_trap_vector(624) <= '1' when (RIN.X.DATA ( 0 ) ( 31 ) /= R_X_DATA031_intermed_1) else '0';
dfp_trap_vector(625) <= '1' when (RIN.X.DATA ( 0 ) ( 31 ) /= R_X_DATA031_intermed_1) else '0';
dfp_trap_vector(626) <= '1' when (RIN.X.DATA ( 0 ) ( 31 ) /= V_X_DATA031_shadow) else '0';
dfp_trap_vector(627) <= '1' when (RIN.X.DATA ( 0 )( 31 ) /= V_X_DATA031_shadow) else '0';
dfp_trap_vector(628) <= '1' when (RIN.X.DATA ( 0 )( 31 ) /= V_X_DATA031_shadow_intermed_1) else '0';
dfp_trap_vector(629) <= '1' when (RIN.X.DATA ( 0 )( 31 ) /= RIN_X_DATA031_intermed_2) else '0';
dfp_trap_vector(630) <= '1' when (RIN.X.DATA ( 0 )( 31 ) /= DCO.DATA ( 0 )( 31 )) else '0';
dfp_trap_vector(631) <= '1' when (RIN.X.DATA ( 0 )( 31 ) /= R_X_DATA031_intermed_1) else '0';
dfp_trap_vector(632) <= '1' when (RIN.X.DATA ( 0 )( 31 ) /= R.X.DATA ( 0 )( 31 )) else '0';
dfp_trap_vector(633) <= '1' when (RIN.E.CTRL.INST ( 19 ) /= DE_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(634) <= '1' when (RIN.E.CTRL.INST ( 19 ) /= V_A_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(635) <= '1' when (RIN.E.CTRL.INST ( 19 ) /= V_E_CTRL_INST19_shadow) else '0';
dfp_trap_vector(636) <= '1' when (RIN.E.CTRL.INST ( 19 ) /= V_E_CTRL_INST19_shadow_intermed_1) else '0';
dfp_trap_vector(637) <= '1' when (RIN.E.CTRL.INST ( 19 ) /= R_E_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(638) <= '1' when (RIN.E.CTRL.INST ( 19 ) /= RIN_A_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(639) <= '1' when (RIN.E.CTRL.INST ( 19 ) /= R_A_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(640) <= '1' when (RIN.E.CTRL.INST ( 19 ) /= R.A.CTRL.INST ( 19 )) else '0';
dfp_trap_vector(641) <= '1' when (RIN.E.CTRL.INST ( 19 ) /= RIN_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(642) <= '1' when (RIN.E.CTRL.INST ( 19 ) /= R.E.CTRL.INST ( 19 )) else '0';
dfp_trap_vector(643) <= '1' when (RIN.E.CTRL.INST ( 19 ) /= RIN_E_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(644) <= '1' when (RIN.E.CTRL.INST ( 19 ) /= V_A_CTRL_INST19_shadow_intermed_1) else '0';
dfp_trap_vector(645) <= '1' when (RIN.E.CTRL.INST ( 20 ) /= V_A_CTRL_INST20_shadow_intermed_1) else '0';
dfp_trap_vector(646) <= '1' when (RIN.E.CTRL.INST ( 20 ) /= R.E.CTRL.INST ( 20 )) else '0';
dfp_trap_vector(647) <= '1' when (RIN.E.CTRL.INST ( 20 ) /= RIN_A_CTRL_INST20_intermed_1) else '0';
dfp_trap_vector(648) <= '1' when (RIN.E.CTRL.INST ( 20 ) /= R.A.CTRL.INST ( 20 )) else '0';
dfp_trap_vector(649) <= '1' when (RIN.E.CTRL.INST ( 20 ) /= R_E_CTRL_INST20_intermed_1) else '0';
dfp_trap_vector(650) <= '1' when (RIN.E.CTRL.INST ( 20 ) /= RIN_A_CTRL_INST20_intermed_2) else '0';
dfp_trap_vector(651) <= '1' when (RIN.E.CTRL.INST ( 20 ) /= V_E_CTRL_INST20_shadow_intermed_1) else '0';
dfp_trap_vector(652) <= '1' when (RIN.E.CTRL.INST ( 20 ) /= V_E_CTRL_INST20_shadow) else '0';
dfp_trap_vector(653) <= '1' when (RIN.E.CTRL.INST ( 20 ) /= DE_INST20_shadow_intermed_2) else '0';
dfp_trap_vector(654) <= '1' when (RIN.E.CTRL.INST ( 20 ) /= V_A_CTRL_INST20_shadow_intermed_2) else '0';
dfp_trap_vector(655) <= '1' when (RIN.E.CTRL.INST ( 20 ) /= RIN_E_CTRL_INST20_intermed_2) else '0';
dfp_trap_vector(656) <= '1' when (RIN.E.CTRL.INST ( 20 ) /= R_A_CTRL_INST20_intermed_1) else '0';
dfp_trap_vector(657) <= '1' when (RIN.X.DATA ( 0 ) ( 0 ) /= RIN_X_DATA00_intermed_2) else '0';
dfp_trap_vector(658) <= '1' when (RIN.X.DATA ( 0 ) ( 0 ) /= V_X_DATA00_shadow) else '0';
dfp_trap_vector(659) <= '1' when (RIN.X.DATA ( 0 ) ( 0 ) /= DCO_DATA00_intermed_1) else '0';
dfp_trap_vector(660) <= '1' when (RIN.X.DATA ( 0 ) ( 0 ) /= V_X_DATA00_shadow_intermed_1) else '0';
dfp_trap_vector(661) <= '1' when (RIN.X.DATA ( 0 ) ( 0 ) /= R.X.DATA ( 0 ) ( 0 )) else '0';
dfp_trap_vector(662) <= '1' when (RIN.X.DATA ( 0 ) ( 0 ) /= V_X_DATA00_shadow_intermed_1) else '0';
dfp_trap_vector(663) <= '1' when (RIN.X.DATA ( 0 ) ( 0 ) /= R_X_DATA00_intermed_1) else '0';
dfp_trap_vector(664) <= '1' when (RIN.X.DATA ( 0 ) ( 0 ) /= RIN_X_DATA00_intermed_2) else '0';
dfp_trap_vector(665) <= '1' when (RIN.X.DATA ( 0 ) ( 0 ) /= R_X_DATA00_intermed_1) else '0';
dfp_trap_vector(666) <= '1' when (RIN.X.DATA ( 0 )( 0 ) /= DCO.DATA ( 0 )( 0 )) else '0';
dfp_trap_vector(667) <= '1' when (RIN.X.DATA ( 0 )( 0 ) /= V_X_DATA00_shadow) else '0';
dfp_trap_vector(668) <= '1' when (RIN.X.DATA ( 0 )( 0 ) /= V_X_DATA00_shadow_intermed_1) else '0';
dfp_trap_vector(669) <= '1' when (RIN.X.DATA ( 0 )( 0 ) /= R.X.DATA ( 0 )( 0 )) else '0';
dfp_trap_vector(670) <= '1' when (RIN.X.DATA ( 0 )( 0 ) /= RIN_X_DATA00_intermed_2) else '0';
dfp_trap_vector(671) <= '1' when (RIN.X.DATA ( 0 )( 0 ) /= R_X_DATA00_intermed_1) else '0';
dfp_trap_vector(672) <= '1' when (RIN.X.DATA ( 0 ) ( 4 DOWNTO 0 ) /= V_X_DATA04DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(673) <= '1' when (RIN.X.DATA ( 0 ) ( 4 DOWNTO 0 ) /= R_X_DATA04DOWNTO0_intermed_1) else '0';
dfp_trap_vector(674) <= '1' when (RIN.X.DATA ( 0 ) ( 4 DOWNTO 0 ) /= R_X_DATA04DOWNTO0_intermed_1) else '0';
dfp_trap_vector(675) <= '1' when (RIN.X.DATA ( 0 ) ( 4 DOWNTO 0 ) /= V_X_DATA04DOWNTO0_shadow) else '0';
dfp_trap_vector(676) <= '1' when (RIN.X.DATA ( 0 ) ( 4 DOWNTO 0 ) /= DCO_DATA04DOWNTO0_intermed_1) else '0';
dfp_trap_vector(677) <= '1' when (RIN.X.DATA ( 0 ) ( 4 DOWNTO 0 ) /= RIN_X_DATA04DOWNTO0_intermed_2) else '0';
dfp_trap_vector(678) <= '1' when (RIN.X.DATA ( 0 ) ( 4 DOWNTO 0 ) /= RIN_X_DATA04DOWNTO0_intermed_2) else '0';
dfp_trap_vector(679) <= '1' when (RIN.X.DATA ( 0 ) ( 4 DOWNTO 0 ) /= R.X.DATA ( 0 ) ( 4 DOWNTO 0 )) else '0';
dfp_trap_vector(680) <= '1' when (RIN.X.DATA ( 0 ) ( 4 DOWNTO 0 ) /= V_X_DATA04DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(681) <= '1' when (RIN.X.DATA ( 0 )( 4 DOWNTO 0 ) /= V_X_DATA04DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(682) <= '1' when (RIN.X.DATA ( 0 )( 4 DOWNTO 0 ) /= R_X_DATA04DOWNTO0_intermed_1) else '0';
dfp_trap_vector(683) <= '1' when (RIN.X.DATA ( 0 )( 4 DOWNTO 0 ) /= R.X.DATA ( 0 )( 4 DOWNTO 0 )) else '0';
dfp_trap_vector(684) <= '1' when (RIN.X.DATA ( 0 )( 4 DOWNTO 0 ) /= DCO.DATA ( 0 )( 4 DOWNTO 0 )) else '0';
dfp_trap_vector(685) <= '1' when (RIN.X.DATA ( 0 )( 4 DOWNTO 0 ) /= RIN_X_DATA04DOWNTO0_intermed_2) else '0';
dfp_trap_vector(686) <= '1' when (RIN.X.DATA ( 0 )( 4 DOWNTO 0 ) /= V_X_DATA04DOWNTO0_shadow) else '0';
dfp_trap_vector(687) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= R_M_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(688) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= RIN_M_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(689) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(690) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= RIN_A_CTRL_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(691) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= R_A_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(692) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(693) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= R_X_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(694) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= V_D_PC31DOWNTO2_shadow_intermed_7) else '0';
dfp_trap_vector(695) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(696) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= RIN_D_PC31DOWNTO2_intermed_7) else '0';
dfp_trap_vector(697) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_1) else '0';
dfp_trap_vector(698) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= V_F_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(699) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= V_F_PC31DOWNTO2_shadow) else '0';
dfp_trap_vector(700) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= RIN_F_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(701) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= RIN_X_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(702) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= IRIN_ADDR31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(703) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= R_E_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(704) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_6) else '0';
dfp_trap_vector(705) <= '1' when (RIN.F.PC ( 2 DOWNTO 2 ) /= "1") else '0';
dfp_trap_vector(706) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(707) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= R_D_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(708) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= R.F.PC ( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(709) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= IR_ADDR31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(710) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= RIN_E_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(711) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= R_F_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(712) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= V_X_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(713) <= '1' when (RIN.F.PC ( 31 DOWNTO 2 ) /= VIR_ADDR31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(714) <= '1' when (RIN.D.PC ( 31 DOWNTO 2 ) /= V_D_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(715) <= '1' when (RIN.D.PC ( 31 DOWNTO 2 ) /= RIN_D_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(716) <= '1' when (RIN.D.PC ( 31 DOWNTO 2 ) /= R.D.PC ( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(717) <= '1' when (RIN.D.PC ( 31 DOWNTO 2 ) /= R_D_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(718) <= '1' when (RIN.D.PC ( 31 DOWNTO 2 ) /= V_D_PC31DOWNTO2_shadow) else '0';
dfp_trap_vector(719) <= '1' when (RIN.E.CTRL.INST ( 24 ) /= V_A_CTRL_INST24_shadow_intermed_2) else '0';
dfp_trap_vector(720) <= '1' when (RIN.E.CTRL.INST ( 24 ) /= V_E_CTRL_INST24_shadow_intermed_1) else '0';
dfp_trap_vector(721) <= '1' when (RIN.E.CTRL.INST ( 24 ) /= DE_INST24_shadow_intermed_2) else '0';
dfp_trap_vector(722) <= '1' when (RIN.E.CTRL.INST ( 24 ) /= V_E_CTRL_INST24_shadow) else '0';
dfp_trap_vector(723) <= '1' when (RIN.E.CTRL.INST ( 24 ) /= R_A_CTRL_INST24_intermed_1) else '0';
dfp_trap_vector(724) <= '1' when (RIN.E.CTRL.INST ( 24 ) /= RIN_A_CTRL_INST24_intermed_1) else '0';
dfp_trap_vector(725) <= '1' when (RIN.E.CTRL.INST ( 24 ) /= V_A_CTRL_INST24_shadow_intermed_1) else '0';
dfp_trap_vector(726) <= '1' when (RIN.E.CTRL.INST ( 24 ) /= RIN_A_CTRL_INST24_intermed_2) else '0';
dfp_trap_vector(727) <= '1' when (RIN.E.CTRL.INST ( 24 ) /= RIN_E_CTRL_INST24_intermed_2) else '0';
dfp_trap_vector(728) <= '1' when (RIN.E.CTRL.INST ( 24 ) /= R_E_CTRL_INST24_intermed_1) else '0';
dfp_trap_vector(729) <= '1' when (RIN.E.CTRL.INST ( 24 ) /= R.A.CTRL.INST ( 24 )) else '0';
dfp_trap_vector(730) <= '1' when (RIN.E.CTRL.INST ( 24 ) /= R.E.CTRL.INST ( 24 )) else '0';
dfp_trap_vector(731) <= '1' when (RIN.A.CTRL.INST ( 19 ) /= DE_INST19_shadow_intermed_1) else '0';
dfp_trap_vector(732) <= '1' when (RIN.A.CTRL.INST ( 19 ) /= V_A_CTRL_INST19_shadow_intermed_1) else '0';
dfp_trap_vector(733) <= '1' when (RIN.A.CTRL.INST ( 19 ) /= R_A_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(734) <= '1' when (RIN.A.CTRL.INST ( 19 ) /= R.A.CTRL.INST ( 19 )) else '0';
dfp_trap_vector(735) <= '1' when (RIN.A.CTRL.INST ( 19 ) /= RIN_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(736) <= '1' when (RIN.A.CTRL.INST ( 19 ) /= V_A_CTRL_INST19_shadow) else '0';
dfp_trap_vector(737) <= '1' when (RIN.M.Y ( 31 ) /= V_M_Y31_shadow_intermed_1) else '0';
dfp_trap_vector(738) <= '1' when (RIN.M.Y ( 31 ) /= V_M_Y31_shadow) else '0';
dfp_trap_vector(739) <= '1' when (RIN.M.Y ( 31 ) /= RIN_M_Y31_intermed_2) else '0';
dfp_trap_vector(740) <= '1' when (RIN.M.Y ( 31 ) /= R_M_Y31_intermed_1) else '0';
dfp_trap_vector(741) <= '1' when (RIN.M.Y ( 31 ) /= R.M.Y ( 31 )) else '0';
dfp_trap_vector(742) <= '1' when (DSUIN.CRDY ( 2 ) /= VDSU_CRDY2_shadow_intermed_1) else '0';
dfp_trap_vector(743) <= '1' when (DSUIN.CRDY ( 2 ) /= VDSU_CRDY2_shadow) else '0';
dfp_trap_vector(744) <= '1' when (DSUIN.CRDY ( 2 ) /= DSUIN_CRDY2_intermed_2) else '0';
dfp_trap_vector(745) <= '1' when (DSUIN.CRDY ( 2 ) /= DSUR.CRDY ( 2 )) else '0';
dfp_trap_vector(746) <= '1' when (DSUIN.CRDY ( 2 ) /= DSUR_CRDY2_intermed_1) else '0';
dfp_trap_vector(747) <= '1' when (RIN.A.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_A_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(748) <= '1' when (RIN.A.CTRL.PC ( 31 DOWNTO 2 ) /= R_A_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(749) <= '1' when (RIN.A.CTRL.PC ( 31 DOWNTO 2 ) /= R.A.CTRL.PC ( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(750) <= '1' when (RIN.A.CTRL.PC ( 31 DOWNTO 2 ) /= V_D_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(751) <= '1' when (RIN.A.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_D_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(752) <= '1' when (RIN.A.CTRL.PC ( 31 DOWNTO 2 ) /= V_A_CTRL_PC31DOWNTO2_shadow) else '0';
dfp_trap_vector(753) <= '1' when (RIN.A.CTRL.PC ( 31 DOWNTO 2 ) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(754) <= '1' when (RIN.A.CTRL.PC ( 31 DOWNTO 2 ) /= R_D_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(755) <= '1' when (RIN.E.CTRL.PC ( 31 DOWNTO 2 ) /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(756) <= '1' when (RIN.E.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_A_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(757) <= '1' when (RIN.E.CTRL.PC ( 31 DOWNTO 2 ) /= R_A_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(758) <= '1' when (RIN.E.CTRL.PC ( 31 DOWNTO 2 ) /= R.A.CTRL.PC ( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(759) <= '1' when (RIN.E.CTRL.PC ( 31 DOWNTO 2 ) /= R.E.CTRL.PC ( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(760) <= '1' when (RIN.E.CTRL.PC ( 31 DOWNTO 2 ) /= V_D_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(761) <= '1' when (RIN.E.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_D_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(762) <= '1' when (RIN.E.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_A_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(763) <= '1' when (RIN.E.CTRL.PC ( 31 DOWNTO 2 ) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(764) <= '1' when (RIN.E.CTRL.PC ( 31 DOWNTO 2 ) /= R_E_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(765) <= '1' when (RIN.E.CTRL.PC ( 31 DOWNTO 2 ) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(766) <= '1' when (RIN.E.CTRL.PC ( 31 DOWNTO 2 ) /= R_D_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(767) <= '1' when (RIN.E.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_E_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(768) <= '1' when (RIN.E.CTRL.PC ( 31 DOWNTO 2 ) /= V_E_CTRL_PC31DOWNTO2_shadow) else '0';
dfp_trap_vector(769) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= R_M_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(770) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_M_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(771) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(772) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_A_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(773) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= V_M_CTRL_PC31DOWNTO2_shadow) else '0';
dfp_trap_vector(774) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= R_A_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(775) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(776) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= R_A_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(777) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= R.E.CTRL.PC ( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(778) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= V_D_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(779) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_D_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(780) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_E_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(781) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_A_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(782) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(783) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= R_E_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(784) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(785) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= R_D_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(786) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= R.M.CTRL.PC ( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(787) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= RIN_E_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(788) <= '1' when (RIN.M.CTRL.PC ( 31 DOWNTO 2 ) /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(789) <= '1' when (R.X.DATA ( 1 ) /= V_X_DATA1_shadow_intermed_1) else '0';
dfp_trap_vector(790) <= '1' when (R.X.DATA ( 1 ) /= DCO_DATA1_intermed_1) else '0';
dfp_trap_vector(791) <= '1' when (R.X.DATA ( 1 ) /= V_X_DATA1_shadow_intermed_2) else '0';
dfp_trap_vector(792) <= '1' when (R.X.DATA ( 1 ) /= RIN_X_DATA1_intermed_1) else '0';
dfp_trap_vector(793) <= '1' when (R.X.DATA ( 1 ) /= R_X_DATA1_intermed_2) else '0';
dfp_trap_vector(794) <= '1' when (R.X.DATA ( 1 ) /= RIN_X_DATA1_intermed_2) else '0';
dfp_trap_vector(795) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= EX_JUMP_ADDRESS31DOWNTO12_shadow_intermed_2) else '0';
dfp_trap_vector(796) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= RIN_F_PC31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(797) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= RIN_A_CTRL_PC31DOWNTO12_intermed_7) else '0';
dfp_trap_vector(798) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= RIN_E_CTRL_PC31DOWNTO12_intermed_6) else '0';
dfp_trap_vector(799) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= V_F_PC31DOWNTO12_shadow_intermed_2) else '0';
dfp_trap_vector(800) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= R_M_CTRL_PC31DOWNTO12_intermed_4) else '0';
dfp_trap_vector(801) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= IRIN_ADDR31DOWNTO12_intermed_3) else '0';
dfp_trap_vector(802) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= V_X_CTRL_PC31DOWNTO12_shadow_intermed_4) else '0';
dfp_trap_vector(803) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= EX_ADD_RES32DOWNTO332DOWNTO13_shadow_intermed_2) else '0';
dfp_trap_vector(804) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= XC_TRAP_ADDRESS31DOWNTO12_shadow_intermed_2) else '0';
dfp_trap_vector(805) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= R_F_PC31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(806) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= RIN_M_CTRL_PC31DOWNTO12_intermed_5) else '0';
dfp_trap_vector(807) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= IR_ADDR31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(808) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= R_X_CTRL_PC31DOWNTO12_intermed_3) else '0';
dfp_trap_vector(809) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= V_D_PC31DOWNTO12_shadow_intermed_8) else '0';
dfp_trap_vector(810) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= V_A_CTRL_PC31DOWNTO12_shadow_intermed_7) else '0';
dfp_trap_vector(811) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= V_E_CTRL_PC31DOWNTO12_shadow_intermed_6) else '0';
dfp_trap_vector(812) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= EX_ADD_RES32DOWNTO330DOWNTO11_shadow_intermed_2) else '0';
dfp_trap_vector(813) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= RIN_F_PC31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(814) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= R_D_PC31DOWNTO12_intermed_7) else '0';
dfp_trap_vector(815) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= R_A_CTRL_PC31DOWNTO12_intermed_6) else '0';
dfp_trap_vector(816) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= R_E_CTRL_PC31DOWNTO12_intermed_5) else '0';
dfp_trap_vector(817) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= RIN_X_CTRL_PC31DOWNTO12_intermed_4) else '0';
dfp_trap_vector(818) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= RIN_D_PC31DOWNTO12_intermed_8) else '0';
dfp_trap_vector(819) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= VIR_ADDR31DOWNTO12_shadow_intermed_3) else '0';
dfp_trap_vector(820) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= V_F_PC31DOWNTO12_shadow_intermed_1) else '0';
dfp_trap_vector(821) <= '1' when (R.F.PC ( 31 DOWNTO 12 ) /= V_M_CTRL_PC31DOWNTO12_shadow_intermed_5) else '0';
dfp_trap_vector(822) <= '1' when (R.D.INST ( 0 ) /= ICO_DATA0_intermed_1) else '0';
dfp_trap_vector(823) <= '1' when (R.D.INST ( 0 ) /= RIN_D_INST0_intermed_1) else '0';
dfp_trap_vector(824) <= '1' when (R.D.INST ( 0 ) /= V_D_INST0_shadow_intermed_2) else '0';
dfp_trap_vector(825) <= '1' when (R.D.INST ( 0 ) /= R_D_INST0_intermed_2) else '0';
dfp_trap_vector(826) <= '1' when (R.D.INST ( 0 ) /= RIN_D_INST0_intermed_2) else '0';
dfp_trap_vector(827) <= '1' when (R.D.INST ( 0 ) /= V_D_INST0_shadow_intermed_1) else '0';
dfp_trap_vector(828) <= '1' when (R.D.INST ( 1 ) /= V_D_INST1_shadow_intermed_2) else '0';
dfp_trap_vector(829) <= '1' when (R.D.INST ( 1 ) /= RIN_D_INST1_intermed_1) else '0';
dfp_trap_vector(830) <= '1' when (R.D.INST ( 1 ) /= RIN_D_INST1_intermed_2) else '0';
dfp_trap_vector(831) <= '1' when (R.D.INST ( 1 ) /= V_D_INST1_shadow_intermed_1) else '0';
dfp_trap_vector(832) <= '1' when (R.D.INST ( 1 ) /= R_D_INST1_intermed_2) else '0';
dfp_trap_vector(833) <= '1' when (R.D.INST ( 1 ) /= ICO_DATA1_intermed_1) else '0';
dfp_trap_vector(834) <= '1' when (R.X.DATA ( 0 )( 31 ) /= RIN_X_DATA031_intermed_1) else '0';
dfp_trap_vector(835) <= '1' when (R.X.DATA ( 0 )( 31 ) /= V_X_DATA031_shadow_intermed_1) else '0';
dfp_trap_vector(836) <= '1' when (R.X.DATA ( 0 )( 31 ) /= V_X_DATA031_shadow_intermed_2) else '0';
dfp_trap_vector(837) <= '1' when (R.X.DATA ( 0 )( 31 ) /= RIN_X_DATA031_intermed_2) else '0';
dfp_trap_vector(838) <= '1' when (R.X.DATA ( 0 )( 31 ) /= DCO_DATA031_intermed_1) else '0';
dfp_trap_vector(839) <= '1' when (R.X.DATA ( 0 )( 31 ) /= R_X_DATA031_intermed_2) else '0';
dfp_trap_vector(840) <= '1' when (RIN.X.DATA ( 1 ) /= V_X_DATA1_shadow) else '0';
dfp_trap_vector(841) <= '1' when (RIN.X.DATA ( 1 ) /= DCO.DATA ( 1 )) else '0';
dfp_trap_vector(842) <= '1' when (RIN.X.DATA ( 1 ) /= V_X_DATA1_shadow_intermed_1) else '0';
dfp_trap_vector(843) <= '1' when (RIN.X.DATA ( 1 ) /= R_X_DATA1_intermed_1) else '0';
dfp_trap_vector(844) <= '1' when (RIN.X.DATA ( 1 ) /= R.X.DATA ( 1 )) else '0';
dfp_trap_vector(845) <= '1' when (RIN.X.DATA ( 1 ) /= RIN_X_DATA1_intermed_2) else '0';
dfp_trap_vector(846) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= EX_JUMP_ADDRESS31DOWNTO12_shadow_intermed_1) else '0';
dfp_trap_vector(847) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= R.F.PC ( 31 DOWNTO 12 )) else '0';
dfp_trap_vector(848) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= RIN_A_CTRL_PC31DOWNTO12_intermed_6) else '0';
dfp_trap_vector(849) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= RIN_E_CTRL_PC31DOWNTO12_intermed_5) else '0';
dfp_trap_vector(850) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= V_F_PC31DOWNTO12_shadow_intermed_1) else '0';
dfp_trap_vector(851) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= R_M_CTRL_PC31DOWNTO12_intermed_3) else '0';
dfp_trap_vector(852) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= IRIN_ADDR31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(853) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= V_X_CTRL_PC31DOWNTO12_shadow_intermed_3) else '0';
dfp_trap_vector(854) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= EX_ADD_RES32DOWNTO332DOWNTO13_shadow_intermed_1) else '0';
dfp_trap_vector(855) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= XC_TRAP_ADDRESS31DOWNTO12_shadow_intermed_1) else '0';
dfp_trap_vector(856) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= R_F_PC31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(857) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= RIN_M_CTRL_PC31DOWNTO12_intermed_4) else '0';
dfp_trap_vector(858) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= IR_ADDR31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(859) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= R_X_CTRL_PC31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(860) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= V_D_PC31DOWNTO12_shadow_intermed_7) else '0';
dfp_trap_vector(861) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= V_A_CTRL_PC31DOWNTO12_shadow_intermed_6) else '0';
dfp_trap_vector(862) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= V_E_CTRL_PC31DOWNTO12_shadow_intermed_5) else '0';
dfp_trap_vector(863) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= EX_ADD_RES32DOWNTO330DOWNTO11_shadow_intermed_1) else '0';
dfp_trap_vector(864) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= RIN_F_PC31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(865) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= R_D_PC31DOWNTO12_intermed_6) else '0';
dfp_trap_vector(866) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= R_A_CTRL_PC31DOWNTO12_intermed_5) else '0';
dfp_trap_vector(867) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= R_E_CTRL_PC31DOWNTO12_intermed_4) else '0';
dfp_trap_vector(868) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= RIN_X_CTRL_PC31DOWNTO12_intermed_3) else '0';
dfp_trap_vector(869) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= RIN_D_PC31DOWNTO12_intermed_7) else '0';
dfp_trap_vector(870) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= VIR_ADDR31DOWNTO12_shadow_intermed_2) else '0';
dfp_trap_vector(871) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= V_F_PC31DOWNTO12_shadow) else '0';
dfp_trap_vector(872) <= '1' when (RIN.F.PC ( 31 DOWNTO 12 ) /= V_M_CTRL_PC31DOWNTO12_shadow_intermed_4) else '0';
dfp_trap_vector(873) <= '1' when (RIN.D.INST ( 0 ) /= ICO.DATA ( 0 )) else '0';
dfp_trap_vector(874) <= '1' when (RIN.D.INST ( 0 ) /= V_D_INST0_shadow_intermed_1) else '0';
dfp_trap_vector(875) <= '1' when (RIN.D.INST ( 0 ) /= R_D_INST0_intermed_1) else '0';
dfp_trap_vector(876) <= '1' when (RIN.D.INST ( 0 ) /= RIN_D_INST0_intermed_2) else '0';
dfp_trap_vector(877) <= '1' when (RIN.D.INST ( 0 ) /= R.D.INST ( 0 )) else '0';
dfp_trap_vector(878) <= '1' when (RIN.D.INST ( 0 ) /= V_D_INST0_shadow) else '0';
dfp_trap_vector(879) <= '1' when (RIN.D.INST ( 1 ) /= V_D_INST1_shadow_intermed_1) else '0';
dfp_trap_vector(880) <= '1' when (RIN.D.INST ( 1 ) /= RIN_D_INST1_intermed_2) else '0';
dfp_trap_vector(881) <= '1' when (RIN.D.INST ( 1 ) /= V_D_INST1_shadow) else '0';
dfp_trap_vector(882) <= '1' when (RIN.D.INST ( 1 ) /= R_D_INST1_intermed_1) else '0';
dfp_trap_vector(883) <= '1' when (RIN.D.INST ( 1 ) /= R.D.INST ( 1 )) else '0';
dfp_trap_vector(884) <= '1' when (RIN.D.INST ( 1 ) /= ICO.DATA ( 1 )) else '0';
dfp_trap_vector(885) <= '1' when (R.X.DATA ( 0 )( 3 ) /= V_X_DATA03_shadow_intermed_2) else '0';
dfp_trap_vector(886) <= '1' when (R.X.DATA ( 0 )( 3 ) /= V_X_DATA03_shadow_intermed_1) else '0';
dfp_trap_vector(887) <= '1' when (R.X.DATA ( 0 )( 3 ) /= DCO_DATA03_intermed_1) else '0';
dfp_trap_vector(888) <= '1' when (R.X.DATA ( 0 )( 3 ) /= RIN_X_DATA03_intermed_1) else '0';
dfp_trap_vector(889) <= '1' when (R.X.DATA ( 0 )( 3 ) /= R_X_DATA03_intermed_2) else '0';
dfp_trap_vector(890) <= '1' when (R.X.DATA ( 0 )( 3 ) /= RIN_X_DATA03_intermed_2) else '0';
dfp_trap_vector(891) <= '1' when (RIN.X.DATA ( 0 )( 3 ) /= V_X_DATA03_shadow_intermed_1) else '0';
dfp_trap_vector(892) <= '1' when (RIN.X.DATA ( 0 )( 3 ) /= V_X_DATA03_shadow) else '0';
dfp_trap_vector(893) <= '1' when (RIN.X.DATA ( 0 )( 3 ) /= DCO.DATA ( 0 )( 3 )) else '0';
dfp_trap_vector(894) <= '1' when (RIN.X.DATA ( 0 )( 3 ) /= R.X.DATA ( 0 )( 3 )) else '0';
dfp_trap_vector(895) <= '1' when (RIN.X.DATA ( 0 )( 3 ) /= R_X_DATA03_intermed_1) else '0';
dfp_trap_vector(896) <= '1' when (RIN.X.DATA ( 0 )( 3 ) /= RIN_X_DATA03_intermed_2) else '0';
dfp_trap_vector(897) <= '1' when (R.A.CTRL.INST ( 20 ) /= V_A_CTRL_INST20_shadow_intermed_1) else '0';
dfp_trap_vector(898) <= '1' when (R.A.CTRL.INST ( 20 ) /= RIN_A_CTRL_INST20_intermed_1) else '0';
dfp_trap_vector(899) <= '1' when (R.A.CTRL.INST ( 20 ) /= RIN_A_CTRL_INST20_intermed_2) else '0';
dfp_trap_vector(900) <= '1' when (R.A.CTRL.INST ( 20 ) /= DE_INST20_shadow_intermed_2) else '0';
dfp_trap_vector(901) <= '1' when (R.A.CTRL.INST ( 20 ) /= V_A_CTRL_INST20_shadow_intermed_2) else '0';
dfp_trap_vector(902) <= '1' when (R.A.CTRL.INST ( 20 ) /= R_A_CTRL_INST20_intermed_2) else '0';
dfp_trap_vector(903) <= '1' when (R.X.DATA ( 0 )( 0 ) /= RIN_X_DATA00_intermed_1) else '0';
dfp_trap_vector(904) <= '1' when (R.X.DATA ( 0 )( 0 ) /= DCO_DATA00_intermed_1) else '0';
dfp_trap_vector(905) <= '1' when (R.X.DATA ( 0 )( 0 ) /= V_X_DATA00_shadow_intermed_1) else '0';
dfp_trap_vector(906) <= '1' when (R.X.DATA ( 0 )( 0 ) /= V_X_DATA00_shadow_intermed_2) else '0';
dfp_trap_vector(907) <= '1' when (R.X.DATA ( 0 )( 0 ) /= RIN_X_DATA00_intermed_2) else '0';
dfp_trap_vector(908) <= '1' when (R.X.DATA ( 0 )( 0 ) /= R_X_DATA00_intermed_2) else '0';
dfp_trap_vector(909) <= '1' when (R.X.DATA ( 0 )( 4 DOWNTO 0 ) /= V_X_DATA04DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(910) <= '1' when (R.X.DATA ( 0 )( 4 DOWNTO 0 ) /= R_X_DATA04DOWNTO0_intermed_2) else '0';
dfp_trap_vector(911) <= '1' when (R.X.DATA ( 0 )( 4 DOWNTO 0 ) /= DCO_DATA04DOWNTO0_intermed_1) else '0';
dfp_trap_vector(912) <= '1' when (R.X.DATA ( 0 )( 4 DOWNTO 0 ) /= RIN_X_DATA04DOWNTO0_intermed_2) else '0';
dfp_trap_vector(913) <= '1' when (R.X.DATA ( 0 )( 4 DOWNTO 0 ) /= RIN_X_DATA04DOWNTO0_intermed_1) else '0';
dfp_trap_vector(914) <= '1' when (R.X.DATA ( 0 )( 4 DOWNTO 0 ) /= V_X_DATA04DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(915) <= '1' when (R.A.CTRL.INST ( 24 ) /= V_A_CTRL_INST24_shadow_intermed_2) else '0';
dfp_trap_vector(916) <= '1' when (R.A.CTRL.INST ( 24 ) /= DE_INST24_shadow_intermed_2) else '0';
dfp_trap_vector(917) <= '1' when (R.A.CTRL.INST ( 24 ) /= R_A_CTRL_INST24_intermed_2) else '0';
dfp_trap_vector(918) <= '1' when (R.A.CTRL.INST ( 24 ) /= RIN_A_CTRL_INST24_intermed_1) else '0';
dfp_trap_vector(919) <= '1' when (R.A.CTRL.INST ( 24 ) /= V_A_CTRL_INST24_shadow_intermed_1) else '0';
dfp_trap_vector(920) <= '1' when (R.A.CTRL.INST ( 24 ) /= RIN_A_CTRL_INST24_intermed_2) else '0';
dfp_trap_vector(921) <= '1' when (RIN.A.CTRL.INST ( 20 ) /= V_A_CTRL_INST20_shadow) else '0';
dfp_trap_vector(922) <= '1' when (RIN.A.CTRL.INST ( 20 ) /= R.A.CTRL.INST ( 20 )) else '0';
dfp_trap_vector(923) <= '1' when (RIN.A.CTRL.INST ( 20 ) /= RIN_A_CTRL_INST20_intermed_2) else '0';
dfp_trap_vector(924) <= '1' when (RIN.A.CTRL.INST ( 20 ) /= DE_INST20_shadow_intermed_1) else '0';
dfp_trap_vector(925) <= '1' when (RIN.A.CTRL.INST ( 20 ) /= V_A_CTRL_INST20_shadow_intermed_1) else '0';
dfp_trap_vector(926) <= '1' when (RIN.A.CTRL.INST ( 20 ) /= R_A_CTRL_INST20_intermed_1) else '0';
dfp_trap_vector(927) <= '1' when (RIN.A.CTRL.INST ( 24 ) /= V_A_CTRL_INST24_shadow_intermed_1) else '0';
dfp_trap_vector(928) <= '1' when (RIN.A.CTRL.INST ( 24 ) /= DE_INST24_shadow_intermed_1) else '0';
dfp_trap_vector(929) <= '1' when (RIN.A.CTRL.INST ( 24 ) /= R_A_CTRL_INST24_intermed_1) else '0';
dfp_trap_vector(930) <= '1' when (RIN.A.CTRL.INST ( 24 ) /= V_A_CTRL_INST24_shadow) else '0';
dfp_trap_vector(931) <= '1' when (RIN.A.CTRL.INST ( 24 ) /= RIN_A_CTRL_INST24_intermed_2) else '0';
dfp_trap_vector(932) <= '1' when (RIN.A.CTRL.INST ( 24 ) /= R.A.CTRL.INST ( 24 )) else '0';
dfp_trap_vector(933) <= '1' when (R.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 ) /= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(934) <= '1' when (R.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 ) /= R_X_RESULT6DOWNTO03DOWNTO0_intermed_2) else '0';
dfp_trap_vector(935) <= '1' when (R.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 ) /= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2) else '0';
dfp_trap_vector(936) <= '1' when (R.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 ) /= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1) else '0';
dfp_trap_vector(937) <= '1' when (R.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 ) /= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(938) <= '1' when (RIN.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 ) /= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(939) <= '1' when (RIN.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 ) /= R_X_RESULT6DOWNTO03DOWNTO0_intermed_1) else '0';
dfp_trap_vector(940) <= '1' when (RIN.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 ) /= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2) else '0';
dfp_trap_vector(941) <= '1' when (RIN.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 ) /= R.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 )) else '0';
dfp_trap_vector(942) <= '1' when (RIN.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 ) /= V_X_RESULT6DOWNTO03DOWNTO0_shadow) else '0';
dfp_trap_vector(943) <= '1' when (NPC_shadow /= RIN_F_PC_intermed_1) else '0';
dfp_trap_vector(944) <= '1' when (NPC_shadow /= EX_ADD_RES32DOWNTO3_shadow_intermed_1) else '0';
dfp_trap_vector(945) <= '1' when (NPC_shadow /= XC_TRAP_ADDRESS_shadow_intermed_1) else '0';
dfp_trap_vector(946) <= '1' when (NPC_shadow /= R.F.PC) else '0';
dfp_trap_vector(947) <= '1' when (NPC_shadow /= EX_JUMP_ADDRESS_shadow_intermed_1) else '0';
dfp_trap_vector(948) <= '1' when (NPC_shadow /= "000000000000000000000000000000") else '0';
dfp_trap_vector(949) <= '1' when (NPC_shadow /= V_F_PC_shadow_intermed_1) else '0';
dfp_trap_vector(950) <= '1' when (DE_REN1_shadow /= RIN_A_RFE1_intermed_1) else '0';
dfp_trap_vector(951) <= '1' when (DE_REN1_shadow /= V_A_RFE1_shadow_intermed_1) else '0';
dfp_trap_vector(952) <= '1' when (DE_REN1_shadow /= R.A.RFE1) else '0';
dfp_trap_vector(953) <= '1' when (DE_REN1_shadow /= '1') else '0';
dfp_trap_vector(954) <= '1' when (DE_REN2_shadow /= RIN_A_RFE2_intermed_1) else '0';
dfp_trap_vector(955) <= '1' when (DE_REN2_shadow /= V_A_RFE2_shadow_intermed_1) else '0';
dfp_trap_vector(956) <= '1' when (DE_REN2_shadow /= R.A.RFE2) else '0';
dfp_trap_vector(957) <= '1' when (EX_ADD_RES_shadow(31 downto 0) /= V_X_DATA0_shadow_intermed_2) else '0';
dfp_trap_vector(958) <= '1' when (EX_ADD_RES_shadow(31 downto 0) /= RIN_X_DATA0_intermed_1) else '0';
dfp_trap_vector(959) <= '1' when (EX_ADD_RES_shadow(31 downto 0) /= V_E_OP1_shadow_intermed_1) else '0';
dfp_trap_vector(960) <= '1' when (EX_ADD_RES_shadow(31 downto 0) /= V_E_OP2_shadow_intermed_1) else '0';
dfp_trap_vector(961) <= '1' when (EX_ADD_RES_shadow(31 downto 0) /= RIN_E_OP2_intermed_1) else '0';
dfp_trap_vector(962) <= '1' when (EX_ADD_RES_shadow(31 downto 0) /= RIN_E_OP1_intermed_1) else '0';
dfp_trap_vector(963) <= '1' when (EX_ADD_RES_shadow(31 downto 0) /= V_X_DATA0_shadow_intermed_1) else '0';
dfp_trap_vector(964) <= '1' when (EX_ADD_RES_shadow(31 downto 0) /= EX_OP1_shadow) else '0';
dfp_trap_vector(965) <= '1' when (EX_ADD_RES_shadow(31 downto 0) /= EX_OP2_shadow) else '0';
dfp_trap_vector(966) <= '1' when (EX_ADD_RES_shadow(0) /= V_E_ALUCIN_shadow_intermed_1) else '0';
dfp_trap_vector(967) <= '1' when (EX_ADD_RES_shadow(31 downto 0) /= R_X_DATA0_intermed_1) else '0';
dfp_trap_vector(968) <= '1' when (EX_ADD_RES_shadow(31 downto 0) /= R.X.DATA ( 0 )) else '0';
dfp_trap_vector(969) <= '1' when (EX_ADD_RES_shadow(0) /= R.E.ALUCIN) else '0';
dfp_trap_vector(970) <= '1' when (EX_ADD_RES_shadow(0) /= RIN_E_ALUCIN_intermed_1) else '0';
dfp_trap_vector(971) <= '1' when (EX_ADD_RES_shadow(31 downto 0) /= X"00000001") else '0';
dfp_trap_vector(972) <= '1' when (EX_ADD_RES_shadow(31 downto 0) /= R.E.OP2) else '0';
dfp_trap_vector(973) <= '1' when (EX_ADD_RES_shadow(31 downto 0) /= DCO_DATA0_intermed_1) else '0';
dfp_trap_vector(974) <= '1' when (EX_ADD_RES_shadow(31 downto 0) /= RIN_X_DATA0_intermed_2) else '0';
dfp_trap_vector(975) <= '1' when (EX_ADD_RES_shadow(31 downto 0) /= R.E.OP1) else '0';
dfp_trap_vector(976) <= '1' when (EX_YMSB_shadow /= RIN_X_DATA00_intermed_2) else '0';
dfp_trap_vector(977) <= '1' when (EX_YMSB_shadow /= V_X_DATA00_shadow_intermed_1) else '0';
dfp_trap_vector(978) <= '1' when (EX_YMSB_shadow /= DCO_DATA00_intermed_1) else '0';
dfp_trap_vector(979) <= '1' when (EX_YMSB_shadow /= V_X_DATA00_shadow_intermed_2) else '0';
dfp_trap_vector(980) <= '1' when (EX_YMSB_shadow /= R.X.DATA ( 0 ) ( 0 )) else '0';
dfp_trap_vector(981) <= '1' when (EX_YMSB_shadow /= V_E_YMSB_shadow_intermed_1) else '0';
dfp_trap_vector(982) <= '1' when (EX_YMSB_shadow /= RIN_X_DATA00_intermed_1) else '0';
dfp_trap_vector(983) <= '1' when (EX_YMSB_shadow /= V_X_DATA00_shadow_intermed_3) else '0';
dfp_trap_vector(984) <= '1' when (EX_YMSB_shadow /= R.E.YMSB) else '0';
dfp_trap_vector(985) <= '1' when (EX_YMSB_shadow /= R_X_DATA00_intermed_1) else '0';
dfp_trap_vector(986) <= '1' when (EX_YMSB_shadow /= RIN_X_DATA00_intermed_3) else '0';
dfp_trap_vector(987) <= '1' when (EX_YMSB_shadow /= R_X_DATA00_intermed_2) else '0';
dfp_trap_vector(988) <= '1' when (EX_YMSB_shadow /= RIN_E_YMSB_intermed_1) else '0';
dfp_trap_vector(989) <= '1' when (EX_OP1_shadow /= V_X_DATA0_shadow_intermed_2) else '0';
dfp_trap_vector(990) <= '1' when (EX_OP1_shadow /= RIN_X_DATA0_intermed_1) else '0';
dfp_trap_vector(991) <= '1' when (EX_OP1_shadow /= V_E_OP1_shadow_intermed_1) else '0';
dfp_trap_vector(992) <= '1' when (EX_OP1_shadow /= RIN_E_OP1_intermed_1) else '0';
dfp_trap_vector(993) <= '1' when (EX_OP1_shadow /= V_X_DATA0_shadow_intermed_1) else '0';
dfp_trap_vector(994) <= '1' when (EX_OP1_shadow /= R_X_DATA0_intermed_1) else '0';
dfp_trap_vector(995) <= '1' when (EX_OP1_shadow /= R.X.DATA ( 0 )) else '0';
dfp_trap_vector(996) <= '1' when (EX_OP1_shadow /= DCO_DATA0_intermed_1) else '0';
dfp_trap_vector(997) <= '1' when (EX_OP1_shadow /= RIN_X_DATA0_intermed_2) else '0';
dfp_trap_vector(998) <= '1' when (EX_OP1_shadow /= R.E.OP1) else '0';
dfp_trap_vector(999) <= '1' when (EX_OP2_shadow /= V_X_DATA0_shadow_intermed_2) else '0';
dfp_trap_vector(1000) <= '1' when (EX_OP2_shadow /= RIN_X_DATA0_intermed_1) else '0';
dfp_trap_vector(1001) <= '1' when (EX_OP2_shadow /= V_E_OP2_shadow_intermed_1) else '0';
dfp_trap_vector(1002) <= '1' when (EX_OP2_shadow /= RIN_E_OP2_intermed_1) else '0';
dfp_trap_vector(1003) <= '1' when (EX_OP2_shadow /= V_X_DATA0_shadow_intermed_1) else '0';
dfp_trap_vector(1004) <= '1' when (EX_OP2_shadow /= R_X_DATA0_intermed_1) else '0';
dfp_trap_vector(1005) <= '1' when (EX_OP2_shadow /= R.X.DATA ( 0 )) else '0';
dfp_trap_vector(1006) <= '1' when (EX_OP2_shadow /= R.E.OP2) else '0';
dfp_trap_vector(1007) <= '1' when (EX_OP2_shadow /= DCO_DATA0_intermed_1) else '0';
dfp_trap_vector(1008) <= '1' when (EX_OP2_shadow /= RIN_X_DATA0_intermed_2) else '0';
dfp_trap_vector(1009) <= '1' when (EX_SHCNT_shadow /= RIN_X_DATA04DOWNTO0_intermed_1) else '0';
dfp_trap_vector(1010) <= '1' when (EX_SHCNT_shadow /= V_X_DATA04DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(1011) <= '1' when (EX_SHCNT_shadow /= R.E.SHCNT) else '0';
dfp_trap_vector(1012) <= '1' when (EX_SHCNT_shadow /= R_X_DATA04DOWNTO0_intermed_2) else '0';
dfp_trap_vector(1013) <= '1' when (EX_SHCNT_shadow /= V_E_SHCNT_shadow_intermed_1) else '0';
dfp_trap_vector(1014) <= '1' when (EX_SHCNT_shadow /= R_X_DATA04DOWNTO0_intermed_1) else '0';
dfp_trap_vector(1015) <= '1' when (EX_SHCNT_shadow /= V_X_DATA04DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(1016) <= '1' when (EX_SHCNT_shadow /= RIN_X_DATA04DOWNTO0_intermed_3) else '0';
dfp_trap_vector(1017) <= '1' when (EX_SHCNT_shadow /= RIN_X_DATA04DOWNTO0_intermed_2) else '0';
dfp_trap_vector(1018) <= '1' when (EX_SHCNT_shadow /= DCO_DATA04DOWNTO0_intermed_1) else '0';
dfp_trap_vector(1019) <= '1' when (EX_SHCNT_shadow /= RIN_E_SHCNT_intermed_1) else '0';
dfp_trap_vector(1020) <= '1' when (EX_SHCNT_shadow /= R.X.DATA ( 0 ) ( 4 DOWNTO 0 )) else '0';
dfp_trap_vector(1021) <= '1' when (EX_SHCNT_shadow /= V_X_DATA04DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(1022) <= '1' when (EX_SARI_shadow /= RIN_X_DATA031_intermed_2) else '0';
dfp_trap_vector(1023) <= '1' when (EX_SARI_shadow /= DE_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(1024) <= '1' when (EX_SARI_shadow /= V_A_CTRL_INST20_shadow_intermed_2) else '0';
dfp_trap_vector(1025) <= '1' when (EX_SARI_shadow /= V_A_CTRL_INST19_shadow_intermed_3) else '0';
dfp_trap_vector(1026) <= '1' when (EX_SARI_shadow /= R.E.CTRL.INST ( 20 )) else '0';
dfp_trap_vector(1027) <= '1' when (EX_SARI_shadow /= RIN_A_CTRL_INST20_intermed_2) else '0';
dfp_trap_vector(1028) <= '1' when (EX_SARI_shadow /= V_X_DATA031_shadow_intermed_2) else '0';
dfp_trap_vector(1029) <= '1' when (EX_SARI_shadow /= V_E_CTRL_INST19_shadow_intermed_1) else '0';
dfp_trap_vector(1030) <= '1' when (EX_SARI_shadow /= V_X_DATA031_shadow_intermed_3) else '0';
dfp_trap_vector(1031) <= '1' when (EX_SARI_shadow /= R.X.DATA ( 0 ) ( 31 )) else '0';
dfp_trap_vector(1032) <= '1' when (EX_SARI_shadow /= V_E_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(1033) <= '1' when (EX_SARI_shadow /= RIN_X_DATA031_intermed_3) else '0';
dfp_trap_vector(1034) <= '1' when (EX_SARI_shadow /= RIN_X_DATA031_intermed_1) else '0';
dfp_trap_vector(1035) <= '1' when (EX_SARI_shadow /= V_E_SARI_shadow_intermed_1) else '0';
dfp_trap_vector(1036) <= '1' when (EX_SARI_shadow /= R_E_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(1037) <= '1' when (EX_SARI_shadow /= DCO_DATA031_intermed_1) else '0';
dfp_trap_vector(1038) <= '1' when (EX_SARI_shadow /= R_X_DATA031_intermed_2) else '0';
dfp_trap_vector(1039) <= '1' when (EX_SARI_shadow /= RIN_E_CTRL_INST20_intermed_1) else '0';
dfp_trap_vector(1040) <= '1' when (EX_SARI_shadow /= RIN_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(1041) <= '1' when (EX_SARI_shadow /= R_E_CTRL_INST20_intermed_1) else '0';
dfp_trap_vector(1042) <= '1' when (EX_SARI_shadow /= R_A_CTRL_INST20_intermed_1) else '0';
dfp_trap_vector(1043) <= '1' when (EX_SARI_shadow /= RIN_A_CTRL_INST20_intermed_3) else '0';
dfp_trap_vector(1044) <= '1' when (EX_SARI_shadow /= R_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(1045) <= '1' when (EX_SARI_shadow /= R.E.SARI) else '0';
dfp_trap_vector(1046) <= '1' when (EX_SARI_shadow /= V_E_CTRL_INST20_shadow_intermed_2) else '0';
dfp_trap_vector(1047) <= '1' when (EX_SARI_shadow /= V_E_CTRL_INST20_shadow_intermed_1) else '0';
dfp_trap_vector(1048) <= '1' when (EX_SARI_shadow /= R_A_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(1049) <= '1' when (EX_SARI_shadow /= DE_INST20_shadow_intermed_2) else '0';
dfp_trap_vector(1050) <= '1' when (EX_SARI_shadow /= RIN_A_CTRL_INST19_intermed_3) else '0';
dfp_trap_vector(1051) <= '1' when (EX_SARI_shadow /= RIN_E_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(1052) <= '1' when (EX_SARI_shadow /= R.E.CTRL.INST ( 19 )) else '0';
dfp_trap_vector(1053) <= '1' when (EX_SARI_shadow /= V_A_CTRL_INST20_shadow_intermed_3) else '0';
dfp_trap_vector(1054) <= '1' when (EX_SARI_shadow /= R_X_DATA031_intermed_1) else '0';
dfp_trap_vector(1055) <= '1' when (EX_SARI_shadow /= RIN_E_SARI_intermed_1) else '0';
dfp_trap_vector(1056) <= '1' when (EX_SARI_shadow /= RIN_E_CTRL_INST20_intermed_2) else '0';
dfp_trap_vector(1057) <= '1' when (EX_SARI_shadow /= V_X_DATA031_shadow_intermed_1) else '0';
dfp_trap_vector(1058) <= '1' when (EX_SARI_shadow /= RIN_E_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(1059) <= '1' when (EX_SARI_shadow /= R_A_CTRL_INST20_intermed_2) else '0';
dfp_trap_vector(1060) <= '1' when (EX_SARI_shadow /= V_A_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(1061) <= '1' when (ME_SIGNED_shadow /= V_M_DCI_SIGNED_shadow_intermed_2) else '0';
dfp_trap_vector(1062) <= '1' when (ME_SIGNED_shadow /= RIN_M_DCI_SIGNED_intermed_2) else '0';
dfp_trap_vector(1063) <= '1' when (ME_SIGNED_shadow /= R_M_DCI_SIGNED_intermed_1) else '0';
dfp_trap_vector(1064) <= '1' when (ME_SIGNED_shadow /= R.X.DCI.SIGNED) else '0';
dfp_trap_vector(1065) <= '1' when (ME_SIGNED_shadow /= V_X_DCI_SIGNED_shadow_intermed_1) else '0';
dfp_trap_vector(1066) <= '1' when (ME_SIGNED_shadow /= RIN_X_DCI_SIGNED_intermed_1) else '0';
dfp_trap_vector(1067) <= '1' when (ME_SIZE_shadow /= R.X.DCI.SIZE) else '0';
dfp_trap_vector(1068) <= '1' when (ME_SIZE_shadow /= RIN_M_DCI_SIZE_intermed_2) else '0';
dfp_trap_vector(1069) <= '1' when (ME_SIZE_shadow /= V_M_DCI_SIZE_shadow_intermed_2) else '0';
dfp_trap_vector(1070) <= '1' when (ME_SIZE_shadow /= R_M_DCI_SIZE_intermed_1) else '0';
dfp_trap_vector(1071) <= '1' when (ME_SIZE_shadow /= V_X_DCI_SIZE_shadow_intermed_1) else '0';
dfp_trap_vector(1072) <= '1' when (ME_SIZE_shadow /= RIN_X_DCI_SIZE_intermed_1) else '0';
dfp_trap_vector(1073) <= '1' when (ME_LADDR_shadow /= V_M_RESULT1DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(1074) <= '1' when (ME_LADDR_shadow /= RIN_X_LADDR_intermed_1) else '0';
dfp_trap_vector(1075) <= '1' when (ME_LADDR_shadow /= R_M_RESULT1DOWNTO0_intermed_1) else '0';
dfp_trap_vector(1076) <= '1' when (ME_LADDR_shadow /= RIN_M_RESULT1DOWNTO0_intermed_2) else '0';
dfp_trap_vector(1077) <= '1' when (ME_LADDR_shadow /= RIN_M_RESULT1DOWNTO0_intermed_3) else '0';
dfp_trap_vector(1078) <= '1' when (ME_LADDR_shadow /= V_M_RESULT1DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(1079) <= '1' when (ME_LADDR_shadow /= V_X_LADDR_shadow_intermed_1) else '0';
dfp_trap_vector(1080) <= '1' when (ME_LADDR_shadow /= R.X.LADDR) else '0';
dfp_trap_vector(1081) <= '1' when (ME_LADDR_shadow /= R_M_RESULT1DOWNTO0_intermed_2) else '0';
dfp_trap_vector(1082) <= '1' when (XC_RESULT_shadow /= V_X_DATA0_shadow_intermed_2) else '0';
dfp_trap_vector(1083) <= '1' when (XC_RESULT_shadow(31 downto 2) /= R_M_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(1084) <= '1' when (XC_RESULT_shadow(31 downto 2) /= RIN_M_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(1085) <= '1' when (XC_RESULT_shadow(31 downto 2) /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(1086) <= '1' when (XC_RESULT_shadow(31 downto 2) /= RIN_A_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(1087) <= '1' when (XC_RESULT_shadow /= RIN_X_RESULT_intermed_1) else '0';
dfp_trap_vector(1088) <= '1' when (XC_RESULT_shadow(31 downto 2) /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(1089) <= '1' when (XC_RESULT_shadow(31 downto 2) /= V_X_CTRL_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(1090) <= '1' when (XC_RESULT_shadow(31 downto 2) /= R_A_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(1091) <= '1' when (XC_RESULT_shadow(31 downto 2) /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(1092) <= '1' when (XC_RESULT_shadow /= RIN_X_DATA0_intermed_1) else '0';
dfp_trap_vector(1093) <= '1' when (XC_RESULT_shadow(31 downto 2) /= R_A_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(1094) <= '1' when (XC_RESULT_shadow /= V_X_RESULT_shadow_intermed_1) else '0';
dfp_trap_vector(1095) <= '1' when (XC_RESULT_shadow(31 downto 2) /= R_X_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(1096) <= '1' when (XC_RESULT_shadow(31 downto 2) /= R_E_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(1097) <= '1' when (XC_RESULT_shadow(31 downto 2) /= V_D_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(1098) <= '1' when (XC_RESULT_shadow(31 downto 2) /= RIN_D_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(1099) <= '1' when (XC_RESULT_shadow /= V_X_DATA0_shadow_intermed_1) else '0';
dfp_trap_vector(1100) <= '1' when (XC_RESULT_shadow /= R.X.RESULT) else '0';
dfp_trap_vector(1101) <= '1' when (XC_RESULT_shadow(31 downto 2) /= RIN_E_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(1102) <= '1' when (XC_RESULT_shadow(31 downto 2) /= RIN_A_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(1103) <= '1' when (XC_RESULT_shadow(31 downto 2) /= RIN_X_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(1104) <= '1' when (XC_RESULT_shadow /= R_X_DATA0_intermed_1) else '0';
dfp_trap_vector(1105) <= '1' when (XC_RESULT_shadow(31 downto 2) /= RIN_X_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(1106) <= '1' when (XC_RESULT_shadow(31 downto 2) /= RIN_M_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(1107) <= '1' when (XC_RESULT_shadow /= R.X.DATA ( 0 )) else '0';
dfp_trap_vector(1108) <= '1' when (XC_RESULT_shadow(31 downto 2) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(1109) <= '1' when (XC_RESULT_shadow /= X"00000000") else '0';
dfp_trap_vector(1110) <= '1' when (XC_RESULT_shadow(31 downto 2) /= R.X.CTRL.PC ( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(1111) <= '1' when (XC_RESULT_shadow(31 downto 2) /= R_E_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(1112) <= '1' when (XC_RESULT_shadow(31 downto 2) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(1113) <= '1' when (XC_RESULT_shadow(31 downto 2) /= R_D_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(1114) <= '1' when (XC_RESULT_shadow(31 downto 2) /= R_M_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(1115) <= '1' when (XC_RESULT_shadow /= DCO_DATA0_intermed_1) else '0';
dfp_trap_vector(1116) <= '1' when (XC_RESULT_shadow(31 downto 2) /= RIN_E_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(1117) <= '1' when (XC_RESULT_shadow(31 downto 2) /= V_X_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(1118) <= '1' when (XC_RESULT_shadow(31 downto 2) /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(1119) <= '1' when (XC_RESULT_shadow /= RIN_X_DATA0_intermed_2) else '0';
dfp_trap_vector(1120) <= '1' when (XC_EXCEPTION_shadow /= '1') else '0';
dfp_trap_vector(1121) <= '1' when (XC_EXCEPTION_shadow /= '0') else '0';
dfp_trap_vector(1122) <= '1' when (XC_WREG_shadow /= V_X_ANNUL_ALL_shadow_intermed_4) else '0';
dfp_trap_vector(1123) <= '1' when (XC_WREG_shadow /= RIN_A_CTRL_ANNUL_intermed_5) else '0';
dfp_trap_vector(1124) <= '1' when (XC_WREG_shadow /= R_M_CTRL_WREG_intermed_1) else '0';
dfp_trap_vector(1125) <= '1' when (XC_WREG_shadow /= R.X.CTRL.WREG) else '0';
dfp_trap_vector(1126) <= '1' when (XC_WREG_shadow /= R_A_CTRL_ANNUL_intermed_4) else '0';
dfp_trap_vector(1127) <= '1' when (XC_WREG_shadow /= RIN_X_ANNUL_ALL_intermed_5) else '0';
dfp_trap_vector(1128) <= '1' when (XC_WREG_shadow /= V_M_CTRL_WREG_shadow_intermed_2) else '0';
dfp_trap_vector(1129) <= '1' when (XC_WREG_shadow /= R_X_ANNUL_ALL_intermed_4) else '0';
dfp_trap_vector(1130) <= '1' when (XC_WREG_shadow /= V_X_CTRL_WREG_shadow_intermed_1) else '0';
dfp_trap_vector(1131) <= '1' when (XC_WREG_shadow /= R_E_CTRL_WREG_intermed_2) else '0';
dfp_trap_vector(1132) <= '1' when (XC_WREG_shadow /= RIN_X_CTRL_WREG_intermed_1) else '0';
dfp_trap_vector(1133) <= '1' when (XC_WREG_shadow /= '1') else '0';
dfp_trap_vector(1134) <= '1' when (XC_WREG_shadow /= '0') else '0';
dfp_trap_vector(1135) <= '1' when (XC_WREG_shadow /= V_A_CTRL_ANNUL_shadow_intermed_4) else '0';
dfp_trap_vector(1136) <= '1' when (XC_WREG_shadow /= RIN_E_CTRL_WREG_intermed_3) else '0';
dfp_trap_vector(1137) <= '1' when (XC_WREG_shadow /= RIN_M_CTRL_WREG_intermed_2) else '0';
dfp_trap_vector(1138) <= '1' when (XC_WREG_shadow /= V_E_CTRL_WREG_shadow_intermed_3) else '0';
dfp_trap_vector(1139) <= '1' when (XC_WREG_shadow /= RIN_A_CTRL_WREG_intermed_4) else '0';
dfp_trap_vector(1140) <= '1' when (XC_WREG_shadow /= V_A_CTRL_WREG_shadow_intermed_4) else '0';
dfp_trap_vector(1141) <= '1' when (XC_WREG_shadow /= R_A_CTRL_WREG_intermed_3) else '0';
dfp_trap_vector(1142) <= '1' when (XC_VECTT_shadow(5 downto 0) /= V_E_CTRL_TT_shadow_intermed_3) else '0';
dfp_trap_vector(1143) <= '1' when (XC_VECTT_shadow(5 downto 0) /= V_X_CTRL_TT_shadow_intermed_1) else '0';
dfp_trap_vector(1144) <= '1' when (XC_VECTT_shadow(6 downto 0) /= V_X_RESULT6DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(1145) <= '1' when (XC_VECTT_shadow(5 downto 0) /= RIN_A_CTRL_TT_intermed_4) else '0';
dfp_trap_vector(1146) <= '1' when (XC_VECTT_shadow(6 downto 0) /= RIN_X_RESULT6DOWNTO0_intermed_2) else '0';
dfp_trap_vector(1147) <= '1' when (XC_VECTT_shadow(5 downto 0) /= RIN_E_CTRL_TT_intermed_3) else '0';
dfp_trap_vector(1148) <= '1' when (XC_VECTT_shadow(5 downto 0) /= V_M_CTRL_TT_shadow_intermed_2) else '0';
dfp_trap_vector(1149) <= '1' when (XC_VECTT_shadow(6 downto 0) /= R_X_RESULT6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(1150) <= '1' when (XC_VECTT_shadow(5 downto 0) /= R_A_CTRL_TT_intermed_3) else '0';
dfp_trap_vector(1151) <= '1' when (XC_VECTT_shadow(5 downto 0) /= V_A_CTRL_TT_shadow_intermed_4) else '0';
dfp_trap_vector(1152) <= '1' when (XC_VECTT_shadow(5 downto 0) /= R_M_CTRL_TT_intermed_1) else '0';
dfp_trap_vector(1153) <= '1' when (XC_VECTT_shadow(5 downto 0) /= RIN_X_CTRL_TT_intermed_1) else '0';
dfp_trap_vector(1154) <= '1' when (XC_VECTT_shadow(6 downto 0) /= RIN_X_RESULT6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(1155) <= '1' when (XC_VECTT_shadow /= "00000000") else '0';
dfp_trap_vector(1156) <= '1' when (XC_VECTT_shadow /= "00001001") else '0';
dfp_trap_vector(1157) <= '1' when (XC_VECTT_shadow(5 downto 0) /= R_E_CTRL_TT_intermed_2) else '0';
dfp_trap_vector(1158) <= '1' when (XC_VECTT_shadow /= X"00") else '0';
dfp_trap_vector(1159) <= '1' when (XC_VECTT_shadow /= X"01") else '0';
dfp_trap_vector(1160) <= '1' when (XC_VECTT_shadow(5 downto 0) /= R.X.CTRL.TT) else '0';
dfp_trap_vector(1161) <= '1' when (XC_VECTT_shadow(5 downto 0) /= RIN_M_CTRL_TT_intermed_2) else '0';
dfp_trap_vector(1162) <= '1' when (XC_VECTT_shadow(6 downto 0) /= V_X_RESULT6DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(1163) <= '1' when (XC_VECTT_shadow(6 downto 0) /= R.X.RESULT ( 6 DOWNTO 0 )) else '0';
dfp_trap_vector(1164) <= '1' when (XC_TRAP_shadow /= R.X.CTRL.TRAP) else '0';
dfp_trap_vector(1165) <= '1' when (XC_TRAP_shadow /= V_M_CTRL_TRAP_shadow_intermed_2) else '0';
dfp_trap_vector(1166) <= '1' when (XC_TRAP_shadow /= RIN_X_CTRL_TRAP_intermed_1) else '0';
dfp_trap_vector(1167) <= '1' when (XC_TRAP_shadow /= V_X_CTRL_TRAP_shadow_intermed_1) else '0';
dfp_trap_vector(1168) <= '1' when (XC_TRAP_shadow /= V_A_CTRL_TRAP_shadow_intermed_4) else '0';
dfp_trap_vector(1169) <= '1' when (XC_TRAP_shadow /= V_X_MEXC_shadow_intermed_1) else '0';
dfp_trap_vector(1170) <= '1' when (XC_TRAP_shadow /= V_D_MEXC_shadow_intermed_5) else '0';
dfp_trap_vector(1171) <= '1' when (XC_TRAP_shadow /= R_A_CTRL_TRAP_intermed_3) else '0';
dfp_trap_vector(1172) <= '1' when (XC_TRAP_shadow /= RIN_X_MEXC_intermed_1) else '0';
dfp_trap_vector(1173) <= '1' when (XC_TRAP_shadow /= RIN_M_CTRL_TRAP_intermed_2) else '0';
dfp_trap_vector(1174) <= '1' when (XC_TRAP_shadow /= R_M_CTRL_TRAP_intermed_1) else '0';
dfp_trap_vector(1175) <= '1' when (XC_TRAP_shadow /= ICO_MEXC_intermed_5) else '0';
dfp_trap_vector(1176) <= '1' when (XC_TRAP_shadow /= R_E_CTRL_TRAP_intermed_2) else '0';
dfp_trap_vector(1177) <= '1' when (XC_TRAP_shadow /= RIN_A_CTRL_TRAP_intermed_4) else '0';
dfp_trap_vector(1178) <= '1' when (XC_TRAP_shadow /= V_E_CTRL_TRAP_shadow_intermed_3) else '0';
dfp_trap_vector(1179) <= '1' when (XC_TRAP_shadow /= RIN_E_CTRL_TRAP_intermed_3) else '0';
dfp_trap_vector(1180) <= '1' when (XC_TRAP_shadow /= R.X.MEXC) else '0';
dfp_trap_vector(1181) <= '1' when (XC_TRAP_shadow /= RIN_D_MEXC_intermed_5) else '0';
dfp_trap_vector(1182) <= '1' when (XC_TRAP_shadow /= R_D_MEXC_intermed_4) else '0';
dfp_trap_vector(1183) <= '1' when (XC_TRAP_shadow /= DCO_MEXC_intermed_1) else '0';
dfp_trap_vector(1184) <= '1' when (XC_HALT_shadow /= DBGI.HALT) else '0';
dfp_trap_vector(1185) <= '1' when (XC_HALT_shadow /= '0') else '0';
dfp_trap_vector(1186) <= '1' when (DSIGN_shadow /= DE_INST19_shadow_intermed_1) else '0';
dfp_trap_vector(1187) <= '1' when (DSIGN_shadow /= V_A_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(1188) <= '1' when (DSIGN_shadow /= V_E_CTRL_INST19_shadow_intermed_1) else '0';
dfp_trap_vector(1189) <= '1' when (DSIGN_shadow /= V_E_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(1190) <= '1' when (DSIGN_shadow /= R_E_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(1191) <= '1' when (DSIGN_shadow /= RIN_A_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(1192) <= '1' when (DSIGN_shadow /= R_A_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(1193) <= '1' when (DSIGN_shadow /= R.A.CTRL.INST ( 19 )) else '0';
dfp_trap_vector(1194) <= '1' when (DSIGN_shadow /= RIN_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(1195) <= '1' when (DSIGN_shadow /= RIN_E_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(1196) <= '1' when (DSIGN_shadow /= R.E.CTRL.INST ( 19 )) else '0';
dfp_trap_vector(1197) <= '1' when (DSIGN_shadow /= RIN_E_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(1198) <= '1' when (DSIGN_shadow /= V_A_CTRL_INST19_shadow_intermed_1) else '0';
dfp_trap_vector(1199) <= '1' when (SIDLE_shadow /= VP_ERROR_shadow_intermed_1) else '0';
dfp_trap_vector(1200) <= '1' when (SIDLE_shadow /= ICO.IDLE) else '0';
dfp_trap_vector(1201) <= '1' when (SIDLE_shadow /= RPIN_PWD_intermed_1) else '0';
dfp_trap_vector(1202) <= '1' when (SIDLE_shadow /= V_X_DEBUG_shadow_intermed_1) else '0';
dfp_trap_vector(1203) <= '1' when (SIDLE_shadow /= RP.PWD) else '0';
dfp_trap_vector(1204) <= '1' when (SIDLE_shadow /= VP_PWD_shadow_intermed_1) else '0';
dfp_trap_vector(1205) <= '1' when (SIDLE_shadow /= DCO.IDLE) else '0';
dfp_trap_vector(1206) <= '1' when (SIDLE_shadow /= '1') else '0';
dfp_trap_vector(1207) <= '1' when (SIDLE_shadow /= R.X.DEBUG) else '0';
dfp_trap_vector(1208) <= '1' when (SIDLE_shadow /= '0') else '0';
dfp_trap_vector(1209) <= '1' when (SIDLE_shadow /= RPIN_ERROR_intermed_1) else '0';
dfp_trap_vector(1210) <= '1' when (SIDLE_shadow /= RP.ERROR) else '0';
dfp_trap_vector(1211) <= '1' when (SIDLE_shadow /= RIN_X_DEBUG_intermed_1) else '0';
dfp_trap_vector(1212) <= '1' when (ICNT_shadow /= HOLDN) else '0';
dfp_trap_vector(1213) <= '1' when (ICNT_shadow /= '0') else '0';
dfp_trap_vector(1214) <= '1' when (V_X_NERROR_shadow /= VP_ERROR_shadow_intermed_1) else '0';
dfp_trap_vector(1215) <= '1' when (V_X_NERROR_shadow /= R.X.NERROR) else '0';
dfp_trap_vector(1216) <= '1' when (V_X_NERROR_shadow /= RIN_X_NERROR_intermed_1) else '0';
dfp_trap_vector(1217) <= '1' when (V_X_NERROR_shadow /= '1') else '0';
dfp_trap_vector(1218) <= '1' when (V_X_NERROR_shadow /= '0') else '0';
dfp_trap_vector(1219) <= '1' when (V_X_NERROR_shadow /= RPIN_ERROR_intermed_1) else '0';
dfp_trap_vector(1220) <= '1' when (V_X_NERROR_shadow /= RP.ERROR) else '0';
dfp_trap_vector(1221) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= V_F_PC31DOWNTO4_shadow_intermed_1) else '0';
dfp_trap_vector(1222) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(9 downto 4) /= V_X_CTRL_TT_shadow_intermed_1) else '0';
dfp_trap_vector(1223) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(9 downto 4) /= V_E_CTRL_TT_shadow_intermed_3) else '0';
dfp_trap_vector(1224) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= X"0000000") else '0';
dfp_trap_vector(1225) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(9 downto 4) /= RIN_A_CTRL_TT_intermed_4) else '0';
dfp_trap_vector(1226) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= V_X_CTRL_PC31DOWNTO4_shadow_intermed_3) else '0';
dfp_trap_vector(1227) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= IR_ADDR31DOWNTO4_intermed_1) else '0';
dfp_trap_vector(1228) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= R.F.PC( 31 DOWNTO 4 )) else '0';
dfp_trap_vector(1229) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(9 downto 4) /= R_A_CTRL_TT_intermed_3) else '0';
dfp_trap_vector(1230) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(11 downto 4) /= XC_VECTT_shadow) else '0';
dfp_trap_vector(1231) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(9 downto 4) /= R_M_CTRL_TT_intermed_1) else '0';
dfp_trap_vector(1232) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= RIN_F_PC31DOWNTO4_intermed_1) else '0';
dfp_trap_vector(1233) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= VIR_ADDR31DOWNTO4_shadow_intermed_2) else '0';
dfp_trap_vector(1234) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(10 downto 4) /= RIN_X_RESULT6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(1235) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= X"0000000") else '0';
dfp_trap_vector(1236) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(9 downto 4) /= R_E_CTRL_TT_intermed_2) else '0';
dfp_trap_vector(1237) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= R_A_CTRL_PC31DOWNTO4_intermed_5) else '0';
dfp_trap_vector(1238) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= RIN_A_CTRL_PC31DOWNTO4_intermed_6) else '0';
dfp_trap_vector(1239) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= R_D_PC31DOWNTO4_intermed_6) else '0';
dfp_trap_vector(1240) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= RIN_X_CTRL_PC31DOWNTO4_intermed_3) else '0';
dfp_trap_vector(1241) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= EX_ADD_RES32DOWNTO332DOWNTO5_shadow_intermed_1) else '0';
dfp_trap_vector(1242) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= X"0000001") else '0';
dfp_trap_vector(1243) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(9 downto 4) /= R.X.CTRL.TT) else '0';
dfp_trap_vector(1244) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(23 downto 4) /= V_W_S_TBA_shadow_intermed_1) else '0';
dfp_trap_vector(1245) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(9 downto 4) /= RIN_M_CTRL_TT_intermed_2) else '0';
dfp_trap_vector(1246) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= RIN_M_CTRL_PC31DOWNTO4_intermed_4) else '0';
dfp_trap_vector(1247) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= V_E_CTRL_PC31DOWNTO4_shadow_intermed_5) else '0';
dfp_trap_vector(1248) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= V_D_PC31DOWNTO4_shadow_intermed_7) else '0';
dfp_trap_vector(1249) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(10 downto 4) /= V_X_RESULT6DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(1250) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(10 downto 4) /= R.X.RESULT ( 6 DOWNTO 0 )) else '0';
dfp_trap_vector(1251) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= R_X_CTRL_PC31DOWNTO4_intermed_2) else '0';
dfp_trap_vector(1252) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(10 downto 4) /= V_X_RESULT6DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(1253) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(10 downto 4) /= RIN_X_RESULT6DOWNTO0_intermed_2) else '0';
dfp_trap_vector(1254) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(23 downto 4) /= R.W.S.TBA) else '0';
dfp_trap_vector(1255) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(9 downto 4) /= RIN_E_CTRL_TT_intermed_3) else '0';
dfp_trap_vector(1256) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(10 downto 4) /= R_X_RESULT6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(1257) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(9 downto 4) /= V_M_CTRL_TT_shadow_intermed_2) else '0';
dfp_trap_vector(1258) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= IRIN_ADDR31DOWNTO4_intermed_2) else '0';
dfp_trap_vector(1259) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= V_M_CTRL_PC31DOWNTO4_shadow_intermed_4) else '0';
dfp_trap_vector(1260) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(9 downto 4) /= V_A_CTRL_TT_shadow_intermed_4) else '0';
dfp_trap_vector(1261) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= XC_TRAP_ADDRESS31DOWNTO4_shadow_intermed_1) else '0';
dfp_trap_vector(1262) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= R_M_CTRL_PC31DOWNTO4_intermed_3) else '0';
dfp_trap_vector(1263) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(9 downto 4) /= RIN_X_CTRL_TT_intermed_1) else '0';
dfp_trap_vector(1264) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= X"0001001") else '0';
dfp_trap_vector(1265) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= RIN_D_PC31DOWNTO4_intermed_7) else '0';
dfp_trap_vector(1266) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= RIN_E_CTRL_PC31DOWNTO4_intermed_5) else '0';
dfp_trap_vector(1267) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= EX_JUMP_ADDRESS31DOWNTO4_shadow_intermed_1) else '0';
dfp_trap_vector(1268) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow(23 downto 4) /= RIN_W_S_TBA_intermed_1) else '0';
dfp_trap_vector(1269) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= V_A_CTRL_PC31DOWNTO4_shadow_intermed_6) else '0';
dfp_trap_vector(1270) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= X"0000000") else '0';
dfp_trap_vector(1271) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= R_E_CTRL_PC31DOWNTO4_intermed_4) else '0';
dfp_trap_vector(1272) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= R_D_PC3DOWNTO2_intermed_6) else '0';
dfp_trap_vector(1273) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= V_D_PC3DOWNTO2_shadow_intermed_7) else '0';
dfp_trap_vector(1274) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= VIR_ADDR3DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(1275) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= RIN_D_PC3DOWNTO2_intermed_7) else '0';
dfp_trap_vector(1276) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= R_M_CTRL_PC3DOWNTO2_intermed_3) else '0';
dfp_trap_vector(1277) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= R_E_CTRL_PC3DOWNTO2_intermed_4) else '0';
dfp_trap_vector(1278) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= V_E_CTRL_PC3DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(1279) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= RIN_X_CTRL_PC3DOWNTO2_intermed_3) else '0';
dfp_trap_vector(1280) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= R_A_CTRL_PC3DOWNTO2_intermed_5) else '0';
dfp_trap_vector(1281) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= R.F.PC( 3 DOWNTO 2 )) else '0';
dfp_trap_vector(1282) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= V_X_CTRL_PC3DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(1283) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= RIN_M_CTRL_PC3DOWNTO2_intermed_4) else '0';
dfp_trap_vector(1284) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= IRIN_ADDR3DOWNTO2_intermed_2) else '0';
dfp_trap_vector(1285) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= EX_JUMP_ADDRESS3DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(1286) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= EX_ADD_RES32DOWNTO34DOWNTO3_shadow_intermed_1) else '0';
dfp_trap_vector(1287) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= RIN_A_CTRL_PC3DOWNTO2_intermed_6) else '0';
dfp_trap_vector(1288) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= XC_TRAP_ADDRESS3DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(1289) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= V_F_PC3DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(1290) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= V_A_CTRL_PC3DOWNTO2_shadow_intermed_6) else '0';
dfp_trap_vector(1291) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= "00") else '0';
dfp_trap_vector(1292) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= IR_ADDR3DOWNTO2_intermed_1) else '0';
dfp_trap_vector(1293) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= V_M_CTRL_PC3DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(1294) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= R_X_CTRL_PC3DOWNTO2_intermed_2) else '0';
dfp_trap_vector(1295) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= RIN_E_CTRL_PC3DOWNTO2_intermed_5) else '0';
dfp_trap_vector(1296) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= RIN_F_PC3DOWNTO2_intermed_1) else '0';
dfp_trap_vector(1297) <= '1' when (V_X_ANNUL_ALL_shadow /= R.X.ANNUL_ALL) else '0';
dfp_trap_vector(1298) <= '1' when (V_X_ANNUL_ALL_shadow /= '1') else '0';
dfp_trap_vector(1299) <= '1' when (V_X_ANNUL_ALL_shadow /= '0') else '0';
dfp_trap_vector(1300) <= '1' when (V_X_ANNUL_ALL_shadow /= RIN_X_ANNUL_ALL_intermed_1) else '0';
dfp_trap_vector(1301) <= '1' when (V_X_DEBUG_shadow /= '1') else '0';
dfp_trap_vector(1302) <= '1' when (V_X_DEBUG_shadow /= R.X.DEBUG) else '0';
dfp_trap_vector(1303) <= '1' when (V_X_DEBUG_shadow /= '0') else '0';
dfp_trap_vector(1304) <= '1' when (V_X_DEBUG_shadow /= RIN_X_DEBUG_intermed_1) else '0';
dfp_trap_vector(1305) <= '1' when (VIR_ADDR_shadow /= RIN_D_PC_intermed_5) else '0';
dfp_trap_vector(1306) <= '1' when (VIR_ADDR_shadow /= RIN_A_CTRL_PC_intermed_4) else '0';
dfp_trap_vector(1307) <= '1' when (VIR_ADDR_shadow /= R_A_CTRL_PC_intermed_3) else '0';
dfp_trap_vector(1308) <= '1' when (VIR_ADDR_shadow /= V_E_CTRL_PC_shadow_intermed_3) else '0';
dfp_trap_vector(1309) <= '1' when (VIR_ADDR_shadow /= IR.ADDR) else '0';
dfp_trap_vector(1310) <= '1' when (VIR_ADDR_shadow /= R_M_CTRL_PC_intermed_1) else '0';
dfp_trap_vector(1311) <= '1' when (VIR_ADDR_shadow /= R.X.CTRL.PC) else '0';
dfp_trap_vector(1312) <= '1' when (VIR_ADDR_shadow /= R_E_CTRL_PC_intermed_2) else '0';
dfp_trap_vector(1313) <= '1' when (VIR_ADDR_shadow /= RIN_M_CTRL_PC_intermed_2) else '0';
dfp_trap_vector(1314) <= '1' when (VIR_ADDR_shadow /= V_X_CTRL_PC_shadow_intermed_1) else '0';
dfp_trap_vector(1315) <= '1' when (VIR_ADDR_shadow /= V_M_CTRL_PC_shadow_intermed_2) else '0';
dfp_trap_vector(1316) <= '1' when (VIR_ADDR_shadow /= V_A_CTRL_PC_shadow_intermed_4) else '0';
dfp_trap_vector(1317) <= '1' when (VIR_ADDR_shadow /= R_D_PC_intermed_4) else '0';
dfp_trap_vector(1318) <= '1' when (VIR_ADDR_shadow /= RIN_E_CTRL_PC_intermed_3) else '0';
dfp_trap_vector(1319) <= '1' when (VIR_ADDR_shadow /= RIN_X_CTRL_PC_intermed_1) else '0';
dfp_trap_vector(1320) <= '1' when (VIR_ADDR_shadow /= V_D_PC_shadow_intermed_5) else '0';
dfp_trap_vector(1321) <= '1' when (VIR_ADDR_shadow /= IRIN_ADDR_intermed_1) else '0';
dfp_trap_vector(1322) <= '1' when (VDSU_TT_shadow(5 downto 0) /= V_E_CTRL_TT_shadow_intermed_3) else '0';
dfp_trap_vector(1323) <= '1' when (VDSU_TT_shadow(5 downto 0) /= V_X_CTRL_TT_shadow_intermed_1) else '0';
dfp_trap_vector(1324) <= '1' when (VDSU_TT_shadow(5 downto 0) /= RIN_A_CTRL_TT_intermed_4) else '0';
dfp_trap_vector(1325) <= '1' when (VDSU_TT_shadow(5 downto 0) /= R_A_CTRL_TT_intermed_3) else '0';
dfp_trap_vector(1326) <= '1' when (VDSU_TT_shadow /= XC_VECTT_shadow) else '0';
dfp_trap_vector(1327) <= '1' when (VDSU_TT_shadow(5 downto 0) /= R_M_CTRL_TT_intermed_1) else '0';
dfp_trap_vector(1328) <= '1' when (VDSU_TT_shadow(6 downto 0) /= RIN_X_RESULT6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(1329) <= '1' when (VDSU_TT_shadow /= DSUIN_TT_intermed_1) else '0';
dfp_trap_vector(1330) <= '1' when (VDSU_TT_shadow /= X"00") else '0';
dfp_trap_vector(1331) <= '1' when (VDSU_TT_shadow(5 downto 0) /= R_E_CTRL_TT_intermed_2) else '0';
dfp_trap_vector(1332) <= '1' when (VDSU_TT_shadow /= X"01") else '0';
dfp_trap_vector(1333) <= '1' when (VDSU_TT_shadow(5 downto 0) /= R.X.CTRL.TT) else '0';
dfp_trap_vector(1334) <= '1' when (VDSU_TT_shadow(5 downto 0) /= RIN_M_CTRL_TT_intermed_2) else '0';
dfp_trap_vector(1335) <= '1' when (VDSU_TT_shadow(6 downto 0) /= V_X_RESULT6DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(1336) <= '1' when (VDSU_TT_shadow(6 downto 0) /= R.X.RESULT ( 6 DOWNTO 0 )) else '0';
dfp_trap_vector(1337) <= '1' when (VDSU_TT_shadow /= DSUR.TT) else '0';
dfp_trap_vector(1338) <= '1' when (VDSU_TT_shadow(6 downto 0) /= V_X_RESULT6DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(1339) <= '1' when (VDSU_TT_shadow(6 downto 0) /= RIN_X_RESULT6DOWNTO0_intermed_2) else '0';
dfp_trap_vector(1340) <= '1' when (VDSU_TT_shadow(5 downto 0) /= RIN_E_CTRL_TT_intermed_3) else '0';
dfp_trap_vector(1341) <= '1' when (VDSU_TT_shadow(5 downto 0) /= V_M_CTRL_TT_shadow_intermed_2) else '0';
dfp_trap_vector(1342) <= '1' when (VDSU_TT_shadow(6 downto 0) /= R_X_RESULT6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(1343) <= '1' when (VDSU_TT_shadow(5 downto 0) /= V_A_CTRL_TT_shadow_intermed_4) else '0';
dfp_trap_vector(1344) <= '1' when (VDSU_TT_shadow(5 downto 0) /= RIN_X_CTRL_TT_intermed_1) else '0';
dfp_trap_vector(1345) <= '1' when (VDSU_TT_shadow /= "00001001") else '0';
dfp_trap_vector(1346) <= '1' when (VDSU_TT_shadow /= X"00") else '0';
dfp_trap_vector(1347) <= '1' when (VP_PWD_shadow /= RP.PWD) else '0';
dfp_trap_vector(1348) <= '1' when (VP_PWD_shadow /= '1') else '0';
dfp_trap_vector(1349) <= '1' when (VP_PWD_shadow /= '0') else '0';
dfp_trap_vector(1350) <= '1' when (VP_PWD_shadow /= RPIN_PWD_intermed_1) else '0';
dfp_trap_vector(1351) <= '1' when (VIR_PWD_shadow /= '1') else '0';
dfp_trap_vector(1352) <= '1' when (VIR_PWD_shadow /= '0') else '0';
dfp_trap_vector(1353) <= '1' when (VIR_PWD_shadow /= IRIN_PWD_intermed_1) else '0';
dfp_trap_vector(1354) <= '1' when (VIR_PWD_shadow /= IR.PWD) else '0';
dfp_trap_vector(1355) <= '1' when (V_W_S_TT_shadow(5 downto 0) /= V_E_CTRL_TT_shadow_intermed_3) else '0';
dfp_trap_vector(1356) <= '1' when (V_W_S_TT_shadow(5 downto 0) /= V_X_CTRL_TT_shadow_intermed_1) else '0';
dfp_trap_vector(1357) <= '1' when (V_W_S_TT_shadow(5 downto 0) /= RIN_A_CTRL_TT_intermed_4) else '0';
dfp_trap_vector(1358) <= '1' when (V_W_S_TT_shadow(5 downto 0) /= R_A_CTRL_TT_intermed_3) else '0';
dfp_trap_vector(1359) <= '1' when (V_W_S_TT_shadow /= XC_VECTT_shadow) else '0';
dfp_trap_vector(1360) <= '1' when (V_W_S_TT_shadow(5 downto 0) /= R_M_CTRL_TT_intermed_1) else '0';
dfp_trap_vector(1361) <= '1' when (V_W_S_TT_shadow(6 downto 0) /= RIN_X_RESULT6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(1362) <= '1' when (V_W_S_TT_shadow /= "00000000") else '0';
dfp_trap_vector(1363) <= '1' when (V_W_S_TT_shadow(5 downto 0) /= R_E_CTRL_TT_intermed_2) else '0';
dfp_trap_vector(1364) <= '1' when (V_W_S_TT_shadow /= X"01") else '0';
dfp_trap_vector(1365) <= '1' when (V_W_S_TT_shadow(5 downto 0) /= R.X.CTRL.TT) else '0';
dfp_trap_vector(1366) <= '1' when (V_W_S_TT_shadow(5 downto 0) /= RIN_M_CTRL_TT_intermed_2) else '0';
dfp_trap_vector(1367) <= '1' when (V_W_S_TT_shadow(6 downto 0) /= V_X_RESULT6DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(1368) <= '1' when (V_W_S_TT_shadow(6 downto 0) /= R.X.RESULT ( 6 DOWNTO 0 )) else '0';
dfp_trap_vector(1369) <= '1' when (V_W_S_TT_shadow(6 downto 0) /= V_X_RESULT6DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(1370) <= '1' when (V_W_S_TT_shadow /= R.W.S.TT) else '0';
dfp_trap_vector(1371) <= '1' when (V_W_S_TT_shadow(6 downto 0) /= RIN_X_RESULT6DOWNTO0_intermed_2) else '0';
dfp_trap_vector(1372) <= '1' when (V_W_S_TT_shadow(5 downto 0) /= RIN_E_CTRL_TT_intermed_3) else '0';
dfp_trap_vector(1373) <= '1' when (V_W_S_TT_shadow(5 downto 0) /= V_M_CTRL_TT_shadow_intermed_2) else '0';
dfp_trap_vector(1374) <= '1' when (V_W_S_TT_shadow(6 downto 0) /= R_X_RESULT6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(1375) <= '1' when (V_W_S_TT_shadow /= RIN_W_S_TT_intermed_1) else '0';
dfp_trap_vector(1376) <= '1' when (V_W_S_TT_shadow(5 downto 0) /= V_A_CTRL_TT_shadow_intermed_4) else '0';
dfp_trap_vector(1377) <= '1' when (V_W_S_TT_shadow(5 downto 0) /= RIN_X_CTRL_TT_intermed_1) else '0';
dfp_trap_vector(1378) <= '1' when (V_W_S_TT_shadow /= "00001001") else '0';
dfp_trap_vector(1379) <= '1' when (V_W_S_TT_shadow /= X"00") else '0';
dfp_trap_vector(1380) <= '1' when (V_W_S_PS_shadow /= '1') else '0';
dfp_trap_vector(1381) <= '1' when (V_W_S_PS_shadow /= R.W.S.S) else '0';
dfp_trap_vector(1382) <= '1' when (V_W_S_PS_shadow /= RIN_W_S_S_intermed_1) else '0';
dfp_trap_vector(1383) <= '1' when (V_W_S_PS_shadow /= RIN_W_S_PS_intermed_1) else '0';
dfp_trap_vector(1384) <= '1' when (V_W_S_PS_shadow /= R.W.S.PS) else '0';
dfp_trap_vector(1385) <= '1' when (V_W_S_PS_shadow /= V_W_S_S_shadow_intermed_1) else '0';
dfp_trap_vector(1386) <= '1' when (V_W_S_S_shadow /= '1') else '0';
dfp_trap_vector(1387) <= '1' when (V_W_S_S_shadow /= R.W.S.S) else '0';
dfp_trap_vector(1388) <= '1' when (V_W_S_S_shadow /= RIN_W_S_S_intermed_1) else '0';
dfp_trap_vector(1389) <= '1' when (XC_WADDR6DOWNTO0_shadow /= RIN_E_CTRL_RD6DOWNTO0_intermed_3) else '0';
dfp_trap_vector(1390) <= '1' when (XC_WADDR6DOWNTO0_shadow /= RIN_M_CTRL_RD6DOWNTO0_intermed_2) else '0';
dfp_trap_vector(1391) <= '1' when (XC_WADDR6DOWNTO0_shadow /= RIN_X_CTRL_RD6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(1392) <= '1' when (XC_WADDR6DOWNTO0_shadow /= V_X_CTRL_RD6DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(1393) <= '1' when (XC_WADDR6DOWNTO0_shadow(2 downto 0) /= RIN_W_S_CWP_intermed_1) else '0';
dfp_trap_vector(1394) <= '1' when (XC_WADDR6DOWNTO0_shadow /= R.X.CTRL.RD( 6 DOWNTO 0 )) else '0';
dfp_trap_vector(1395) <= '1' when (XC_WADDR6DOWNTO0_shadow /= "0000001") else '0';
dfp_trap_vector(1396) <= '1' when (XC_WADDR6DOWNTO0_shadow /= V_M_CTRL_RD6DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(1397) <= '1' when (XC_WADDR6DOWNTO0_shadow /= "0000001") else '0';
dfp_trap_vector(1398) <= '1' when (XC_WADDR6DOWNTO0_shadow /= R_E_CTRL_RD6DOWNTO0_intermed_2) else '0';
dfp_trap_vector(1399) <= '1' when (XC_WADDR6DOWNTO0_shadow /= "0000010") else '0';
dfp_trap_vector(1400) <= '1' when (XC_WADDR6DOWNTO0_shadow /= V_E_CTRL_RD6DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(1401) <= '1' when (XC_WADDR6DOWNTO0_shadow /= V_A_CTRL_RD6DOWNTO0_shadow_intermed_4) else '0';
dfp_trap_vector(1402) <= '1' when (XC_WADDR6DOWNTO0_shadow /= R_A_CTRL_RD6DOWNTO0_intermed_3) else '0';
dfp_trap_vector(1403) <= '1' when (XC_WADDR6DOWNTO0_shadow(2 downto 0) /= R.W.S.CWP) else '0';
dfp_trap_vector(1404) <= '1' when (XC_WADDR6DOWNTO0_shadow /= RIN_A_CTRL_RD6DOWNTO0_intermed_4) else '0';
dfp_trap_vector(1405) <= '1' when (XC_WADDR6DOWNTO0_shadow /= R_M_CTRL_RD6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(1406) <= '1' when (XC_WADDR6DOWNTO0_shadow(2 downto 0) /= V_W_S_CWP_shadow_intermed_1) else '0';
dfp_trap_vector(1407) <= '1' when (V_W_S_ET_shadow /= '0') else '0';
dfp_trap_vector(1408) <= '1' when (V_W_S_ET_shadow /= RIN_W_S_ET_intermed_1) else '0';
dfp_trap_vector(1409) <= '1' when (V_W_S_ET_shadow /= R.W.S.ET) else '0';
dfp_trap_vector(1410) <= '1' when (V_W_S_CWP_shadow /= RIN_W_S_CWP_intermed_1) else '0';
dfp_trap_vector(1411) <= '1' when (V_W_S_CWP_shadow /= "001") else '0';
dfp_trap_vector(1412) <= '1' when (V_W_S_CWP_shadow /= R.W.S.CWP) else '0';
dfp_trap_vector(1413) <= '1' when (VP_ERROR_shadow /= '1') else '0';
dfp_trap_vector(1414) <= '1' when (VP_ERROR_shadow /= '0') else '0';
dfp_trap_vector(1415) <= '1' when (VP_ERROR_shadow /= RP.ERROR) else '0';
dfp_trap_vector(1416) <= '1' when (VP_ERROR_shadow /= RPIN_ERROR_intermed_1) else '0';
dfp_trap_vector(1417) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= RIN_D_PC_intermed_6) else '0';
dfp_trap_vector(1418) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= RIN_M_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(1419) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= VIR_ADDR_shadow_intermed_1) else '0';
dfp_trap_vector(1420) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= RIN_A_CTRL_PC_intermed_5) else '0';
dfp_trap_vector(1421) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= R_A_CTRL_PC_intermed_4) else '0';
dfp_trap_vector(1422) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= V_D_PC31DOWNTO2_shadow_intermed_7) else '0';
dfp_trap_vector(1423) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= V_E_CTRL_PC_shadow_intermed_4) else '0';
dfp_trap_vector(1424) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= EX_ADD_RES32DOWNTO3_shadow_intermed_1) else '0';
dfp_trap_vector(1425) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= XC_TRAP_ADDRESS_shadow_intermed_1) else '0';
dfp_trap_vector(1426) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= RIN_D_PC31DOWNTO2_intermed_7) else '0';
dfp_trap_vector(1427) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_1) else '0';
dfp_trap_vector(1428) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= IR.ADDR) else '0';
dfp_trap_vector(1429) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= V_F_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(1430) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= RIN_F_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(1431) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= R_M_CTRL_PC_intermed_2) else '0';
dfp_trap_vector(1432) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= RIN_X_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(1433) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= R_X_CTRL_PC_intermed_1) else '0';
dfp_trap_vector(1434) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= R_E_CTRL_PC_intermed_3) else '0';
dfp_trap_vector(1435) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= IRIN_ADDR31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(1436) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_6) else '0';
dfp_trap_vector(1437) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= RIN_M_CTRL_PC_intermed_3) else '0';
dfp_trap_vector(1438) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= R_D_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(1439) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= R.F.PC( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(1440) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= VIR_ADDR31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(1441) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= V_X_CTRL_PC_shadow_intermed_2) else '0';
dfp_trap_vector(1442) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= R_M_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(1443) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(1444) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= RIN_A_CTRL_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(1445) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= R_A_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(1446) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= V_M_CTRL_PC_shadow_intermed_3) else '0';
dfp_trap_vector(1447) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(1448) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= V_A_CTRL_PC_shadow_intermed_5) else '0';
dfp_trap_vector(1449) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= R_X_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(1450) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= R_D_PC_intermed_5) else '0';
dfp_trap_vector(1451) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= RIN_F_PC_intermed_1) else '0';
dfp_trap_vector(1452) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(1453) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= RIN_E_CTRL_PC_intermed_4) else '0';
dfp_trap_vector(1454) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= RIN_X_CTRL_PC_intermed_2) else '0';
dfp_trap_vector(1455) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= R.F.PC) else '0';
dfp_trap_vector(1456) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= V_D_PC_shadow_intermed_6) else '0';
dfp_trap_vector(1457) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= R_E_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(1458) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= IRIN_ADDR_intermed_1) else '0';
dfp_trap_vector(1459) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= EX_JUMP_ADDRESS_shadow_intermed_1) else '0';
dfp_trap_vector(1460) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= "000000000000000000000000000000") else '0';
dfp_trap_vector(1461) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(1462) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= IR_ADDR31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(1463) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= V_F_PC_shadow_intermed_1) else '0';
dfp_trap_vector(1464) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= RIN_E_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(1465) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= V_X_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(1466) <= '1' when (VDSU_TBUFCNT_shadow /= DSUR.TBUFCNT) else '0';
dfp_trap_vector(1467) <= '1' when (VDSU_TBUFCNT_shadow /= TBUFCNTX_shadow) else '0';
dfp_trap_vector(1468) <= '1' when (VDSU_TBUFCNT_shadow /= DSUIN_TBUFCNT_intermed_1) else '0';
dfp_trap_vector(1469) <= '1' when (V_W_EXCEPT_shadow /= R.W.EXCEPT) else '0';
dfp_trap_vector(1470) <= '1' when (V_W_EXCEPT_shadow /= XC_EXCEPTION_shadow) else '0';
dfp_trap_vector(1471) <= '1' when (V_W_EXCEPT_shadow /= '1') else '0';
dfp_trap_vector(1472) <= '1' when (V_W_EXCEPT_shadow /= RIN_W_EXCEPT_intermed_1) else '0';
dfp_trap_vector(1473) <= '1' when (V_W_EXCEPT_shadow /= '0') else '0';
dfp_trap_vector(1474) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= RIN_M_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(1475) <= '1' when (V_W_RESULT_shadow /= RIN_X_RESULT_intermed_1) else '0';
dfp_trap_vector(1476) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(1477) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= V_X_CTRL_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(1478) <= '1' when (V_W_RESULT_shadow /= R.W.RESULT) else '0';
dfp_trap_vector(1479) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= R_E_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(1480) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= V_D_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(1481) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= RIN_D_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(1482) <= '1' when (V_W_RESULT_shadow /= V_X_DATA0_shadow_intermed_1) else '0';
dfp_trap_vector(1483) <= '1' when (V_W_RESULT_shadow /= R.X.RESULT) else '0';
dfp_trap_vector(1484) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= RIN_E_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(1485) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= RIN_A_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(1486) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= RIN_X_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(1487) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= RIN_X_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(1488) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= RIN_M_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(1489) <= '1' when (V_W_RESULT_shadow /= R.X.DATA ( 0 )) else '0';
dfp_trap_vector(1490) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= R.X.CTRL.PC ( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(1491) <= '1' when (V_W_RESULT_shadow /= XC_RESULT_shadow) else '0';
dfp_trap_vector(1492) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(1493) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= R_D_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(1494) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= R_M_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(1495) <= '1' when (V_W_RESULT_shadow /= DCO_DATA0_intermed_1) else '0';
dfp_trap_vector(1496) <= '1' when (V_W_RESULT_shadow /= V_X_DATA0_shadow_intermed_2) else '0';
dfp_trap_vector(1497) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= R_M_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(1498) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(1499) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= RIN_A_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(1500) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= R_A_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(1501) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(1502) <= '1' when (V_W_RESULT_shadow /= RIN_X_DATA0_intermed_1) else '0';
dfp_trap_vector(1503) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= R_A_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(1504) <= '1' when (V_W_RESULT_shadow /= V_X_RESULT_shadow_intermed_1) else '0';
dfp_trap_vector(1505) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= R_X_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(1506) <= '1' when (V_W_RESULT_shadow /= RIN_W_RESULT_intermed_1) else '0';
dfp_trap_vector(1507) <= '1' when (V_W_RESULT_shadow /= R_X_DATA0_intermed_1) else '0';
dfp_trap_vector(1508) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(1509) <= '1' when (V_W_RESULT_shadow /= X"00000000") else '0';
dfp_trap_vector(1510) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= R_E_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(1511) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= RIN_E_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(1512) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= V_X_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(1513) <= '1' when (V_W_RESULT_shadow(31 downto 2) /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(1514) <= '1' when (V_W_RESULT_shadow /= RIN_X_DATA0_intermed_2) else '0';
dfp_trap_vector(1515) <= '1' when (V_W_WA_shadow /= V_M_CTRL_RD7DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(1516) <= '1' when (V_W_WA_shadow /= V_E_CTRL_RD7DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(1517) <= '1' when (V_W_WA_shadow /= R_E_CTRL_RD7DOWNTO0_intermed_2) else '0';
dfp_trap_vector(1518) <= '1' when (V_W_WA_shadow /= V_X_CTRL_RD7DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(1519) <= '1' when (V_W_WA_shadow /= R.X.CTRL.RD ( 7 DOWNTO 0 )) else '0';
dfp_trap_vector(1520) <= '1' when (V_W_WA_shadow /= V_A_CTRL_RD7DOWNTO0_shadow_intermed_4) else '0';
dfp_trap_vector(1521) <= '1' when (V_W_WA_shadow /= RIN_W_WA_intermed_1) else '0';
dfp_trap_vector(1522) <= '1' when (V_W_WA_shadow /= RIN_A_CTRL_RD7DOWNTO0_intermed_4) else '0';
dfp_trap_vector(1523) <= '1' when (V_W_WA_shadow /= R_M_CTRL_RD7DOWNTO0_intermed_1) else '0';
dfp_trap_vector(1524) <= '1' when (V_W_WA_shadow /= R_A_CTRL_RD7DOWNTO0_intermed_3) else '0';
dfp_trap_vector(1525) <= '1' when (V_W_WA_shadow /= RIN_E_CTRL_RD7DOWNTO0_intermed_3) else '0';
dfp_trap_vector(1526) <= '1' when (V_W_WA_shadow /= RIN_X_CTRL_RD7DOWNTO0_intermed_1) else '0';
dfp_trap_vector(1527) <= '1' when (V_W_WA_shadow /= RIN_M_CTRL_RD7DOWNTO0_intermed_2) else '0';
dfp_trap_vector(1528) <= '1' when (V_W_WA_shadow /= R.W.WA) else '0';
dfp_trap_vector(1529) <= '1' when (V_W_WA_shadow /= XC_WADDR7DOWNTO0_shadow) else '0';
dfp_trap_vector(1530) <= '1' when (V_W_WREG_shadow /= RIN_A_CTRL_ANNUL_intermed_5) else '0';
dfp_trap_vector(1531) <= '1' when (V_W_WREG_shadow /= R.X.CTRL.WREG) else '0';
dfp_trap_vector(1532) <= '1' when (V_W_WREG_shadow /= R_A_CTRL_ANNUL_intermed_4) else '0';
dfp_trap_vector(1533) <= '1' when (V_W_WREG_shadow /= R.W.WREG) else '0';
dfp_trap_vector(1534) <= '1' when (V_W_WREG_shadow /= R_X_ANNUL_ALL_intermed_4) else '0';
dfp_trap_vector(1535) <= '1' when (V_W_WREG_shadow /= V_X_CTRL_WREG_shadow_intermed_1) else '0';
dfp_trap_vector(1536) <= '1' when (V_W_WREG_shadow /= RIN_X_CTRL_WREG_intermed_1) else '0';
dfp_trap_vector(1537) <= '1' when (V_W_WREG_shadow /= '1') else '0';
dfp_trap_vector(1538) <= '1' when (V_W_WREG_shadow /= '0') else '0';
dfp_trap_vector(1539) <= '1' when (V_W_WREG_shadow /= XC_WREG_shadow) else '0';
dfp_trap_vector(1540) <= '1' when (V_W_WREG_shadow /= RIN_M_CTRL_WREG_intermed_2) else '0';
dfp_trap_vector(1541) <= '1' when (V_W_WREG_shadow /= RIN_A_CTRL_WREG_intermed_4) else '0';
dfp_trap_vector(1542) <= '1' when (V_W_WREG_shadow /= V_A_CTRL_WREG_shadow_intermed_4) else '0';
dfp_trap_vector(1543) <= '1' when (V_W_WREG_shadow /= R_A_CTRL_WREG_intermed_3) else '0';
dfp_trap_vector(1544) <= '1' when (V_W_WREG_shadow /= RIN_W_WREG_intermed_1) else '0';
dfp_trap_vector(1545) <= '1' when (V_W_WREG_shadow /= V_X_ANNUL_ALL_shadow_intermed_4) else '0';
dfp_trap_vector(1546) <= '1' when (V_W_WREG_shadow /= R_M_CTRL_WREG_intermed_1) else '0';
dfp_trap_vector(1547) <= '1' when (V_W_WREG_shadow /= RIN_X_ANNUL_ALL_intermed_5) else '0';
dfp_trap_vector(1548) <= '1' when (V_W_WREG_shadow /= V_M_CTRL_WREG_shadow_intermed_2) else '0';
dfp_trap_vector(1549) <= '1' when (V_W_WREG_shadow /= HOLDN) else '0';
dfp_trap_vector(1550) <= '1' when (V_W_WREG_shadow /= R_E_CTRL_WREG_intermed_2) else '0';
dfp_trap_vector(1551) <= '1' when (V_W_WREG_shadow /= V_A_CTRL_ANNUL_shadow_intermed_4) else '0';
dfp_trap_vector(1552) <= '1' when (V_W_WREG_shadow /= RIN_E_CTRL_WREG_intermed_3) else '0';
dfp_trap_vector(1553) <= '1' when (V_W_WREG_shadow /= V_E_CTRL_WREG_shadow_intermed_3) else '0';
dfp_trap_vector(1554) <= '1' when (V_W_S_SVT_shadow /= R.W.S.SVT) else '0';
dfp_trap_vector(1555) <= '1' when (V_W_S_SVT_shadow /= '0') else '0';
dfp_trap_vector(1556) <= '1' when (V_W_S_SVT_shadow /= RIN_W_S_SVT_intermed_1) else '0';
dfp_trap_vector(1557) <= '1' when (V_W_S_DWT_shadow /= RIN_W_S_DWT_intermed_1) else '0';
dfp_trap_vector(1558) <= '1' when (V_W_S_DWT_shadow /= R.W.S.DWT) else '0';
dfp_trap_vector(1559) <= '1' when (V_W_S_DWT_shadow /= '0') else '0';
dfp_trap_vector(1560) <= '1' when (V_W_S_EF_shadow /= '0') else '0';
dfp_trap_vector(1561) <= '1' when (V_W_S_EF_shadow /= R.W.S.EF) else '0';
dfp_trap_vector(1562) <= '1' when (V_W_S_EF_shadow /= RIN_W_S_EF_intermed_1) else '0';
dfp_trap_vector(1563) <= '1' when (V_X_CTRL_shadow /= RIN_E_CTRL_intermed_2) else '0';
dfp_trap_vector(1564) <= '1' when (V_X_CTRL_shadow /= R_E_CTRL_intermed_1) else '0';
dfp_trap_vector(1565) <= '1' when (V_X_CTRL_shadow /= RIN_X_CTRL_intermed_1) else '0';
dfp_trap_vector(1566) <= '1' when (V_X_CTRL_shadow /= R.M.CTRL) else '0';
dfp_trap_vector(1567) <= '1' when (V_X_CTRL_shadow /= RIN_M_CTRL_intermed_1) else '0';
dfp_trap_vector(1568) <= '1' when (V_X_CTRL_shadow /= V_E_CTRL_shadow_intermed_2) else '0';
dfp_trap_vector(1569) <= '1' when (V_X_CTRL_shadow /= RIN_A_CTRL_intermed_3) else '0';
dfp_trap_vector(1570) <= '1' when (V_X_CTRL_shadow /= R.X.CTRL) else '0';
dfp_trap_vector(1571) <= '1' when (V_X_CTRL_shadow /= V_M_CTRL_shadow_intermed_1) else '0';
dfp_trap_vector(1572) <= '1' when (V_X_CTRL_shadow /= V_A_CTRL_shadow_intermed_3) else '0';
dfp_trap_vector(1573) <= '1' when (V_X_CTRL_shadow /= R_A_CTRL_intermed_2) else '0';
dfp_trap_vector(1574) <= '1' when (V_X_DCI_shadow /= V_M_DCI_shadow_intermed_1) else '0';
dfp_trap_vector(1575) <= '1' when (V_X_DCI_shadow /= RIN_M_DCI_intermed_1) else '0';
dfp_trap_vector(1576) <= '1' when (V_X_DCI_shadow /= RIN_X_DCI_intermed_1) else '0';
dfp_trap_vector(1577) <= '1' when (V_X_DCI_shadow /= R.M.DCI) else '0';
dfp_trap_vector(1578) <= '1' when (V_X_DCI_shadow /= R.X.DCI) else '0';
dfp_trap_vector(1579) <= '1' when (V_X_CTRL_RETT_shadow /= R.M.CTRL.RETT) else '0';
dfp_trap_vector(1580) <= '1' when (V_X_CTRL_RETT_shadow /= RIN_A_CTRL_ANNUL_intermed_4) else '0';
dfp_trap_vector(1581) <= '1' when (V_X_CTRL_RETT_shadow /= R_A_CTRL_ANNUL_intermed_3) else '0';
dfp_trap_vector(1582) <= '1' when (V_X_CTRL_RETT_shadow /= RIN_M_CTRL_RETT_intermed_1) else '0';
dfp_trap_vector(1583) <= '1' when (V_X_CTRL_RETT_shadow /= V_M_CTRL_ANNUL_shadow_intermed_1) else '0';
dfp_trap_vector(1584) <= '1' when (V_X_CTRL_RETT_shadow /= R_X_ANNUL_ALL_intermed_3) else '0';
dfp_trap_vector(1585) <= '1' when (V_X_CTRL_RETT_shadow /= R.M.CTRL.ANNUL) else '0';
dfp_trap_vector(1586) <= '1' when (V_X_CTRL_RETT_shadow /= '1') else '0';
dfp_trap_vector(1587) <= '1' when (V_X_CTRL_RETT_shadow /= '0') else '0';
dfp_trap_vector(1588) <= '1' when (V_X_CTRL_RETT_shadow /= RIN_M_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(1589) <= '1' when (V_X_CTRL_RETT_shadow /= V_E_CTRL_RETT_shadow_intermed_2) else '0';
dfp_trap_vector(1590) <= '1' when (V_X_CTRL_RETT_shadow /= V_A_CTRL_RETT_shadow_intermed_3) else '0';
dfp_trap_vector(1591) <= '1' when (V_X_CTRL_RETT_shadow /= RIN_A_CTRL_RETT_intermed_3) else '0';
dfp_trap_vector(1592) <= '1' when (V_X_CTRL_RETT_shadow /= V_X_ANNUL_ALL_shadow_intermed_3) else '0';
dfp_trap_vector(1593) <= '1' when (V_X_CTRL_RETT_shadow /= RIN_E_CTRL_ANNUL_intermed_2) else '0';
dfp_trap_vector(1594) <= '1' when (V_X_CTRL_RETT_shadow /= R_E_CTRL_RETT_intermed_1) else '0';
dfp_trap_vector(1595) <= '1' when (V_X_CTRL_RETT_shadow /= R.X.CTRL.RETT) else '0';
dfp_trap_vector(1596) <= '1' when (V_X_CTRL_RETT_shadow /= RIN_X_ANNUL_ALL_intermed_4) else '0';
dfp_trap_vector(1597) <= '1' when (V_X_CTRL_RETT_shadow /= RIN_E_CTRL_RETT_intermed_2) else '0';
dfp_trap_vector(1598) <= '1' when (V_X_CTRL_RETT_shadow /= V_E_CTRL_ANNUL_shadow_intermed_2) else '0';
dfp_trap_vector(1599) <= '1' when (V_X_CTRL_RETT_shadow /= V_A_CTRL_ANNUL_shadow_intermed_3) else '0';
dfp_trap_vector(1600) <= '1' when (V_X_CTRL_RETT_shadow /= RIN_X_CTRL_RETT_intermed_1) else '0';
dfp_trap_vector(1601) <= '1' when (V_X_CTRL_RETT_shadow /= V_M_CTRL_RETT_shadow_intermed_1) else '0';
dfp_trap_vector(1602) <= '1' when (V_X_CTRL_RETT_shadow /= R_A_CTRL_RETT_intermed_2) else '0';
dfp_trap_vector(1603) <= '1' when (V_X_CTRL_RETT_shadow /= R_E_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(1604) <= '1' when (V_X_MAC_shadow /= V_E_MAC_shadow_intermed_2) else '0';
dfp_trap_vector(1605) <= '1' when (V_X_MAC_shadow /= RIN_M_MAC_intermed_1) else '0';
dfp_trap_vector(1606) <= '1' when (V_X_MAC_shadow /= RIN_E_MAC_intermed_2) else '0';
dfp_trap_vector(1607) <= '1' when (V_X_MAC_shadow /= R_E_MAC_intermed_1) else '0';
dfp_trap_vector(1608) <= '1' when (V_X_MAC_shadow /= R.M.MAC) else '0';
dfp_trap_vector(1609) <= '1' when (V_X_MAC_shadow /= V_M_MAC_shadow_intermed_1) else '0';
dfp_trap_vector(1610) <= '1' when (V_X_MAC_shadow /= RIN_X_MAC_intermed_1) else '0';
dfp_trap_vector(1611) <= '1' when (V_X_MAC_shadow /= R.X.MAC) else '0';
dfp_trap_vector(1612) <= '1' when (V_X_LADDR_shadow /= V_M_RESULT1DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(1613) <= '1' when (V_X_LADDR_shadow /= RIN_X_LADDR_intermed_1) else '0';
dfp_trap_vector(1614) <= '1' when (V_X_LADDR_shadow /= R.M.RESULT ( 1 DOWNTO 0 )) else '0';
dfp_trap_vector(1615) <= '1' when (V_X_LADDR_shadow /= RIN_M_RESULT1DOWNTO0_intermed_2) else '0';
dfp_trap_vector(1616) <= '1' when (V_X_LADDR_shadow /= V_M_RESULT1DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(1617) <= '1' when (V_X_LADDR_shadow /= R.X.LADDR) else '0';
dfp_trap_vector(1618) <= '1' when (V_X_LADDR_shadow /= R_M_RESULT1DOWNTO0_intermed_1) else '0';
dfp_trap_vector(1619) <= '1' when (V_X_LADDR_shadow /= RIN_M_RESULT1DOWNTO0_intermed_1) else '0';
dfp_trap_vector(1620) <= '1' when (V_X_CTRL_ANNUL_shadow /= RIN_A_CTRL_ANNUL_intermed_3) else '0';
dfp_trap_vector(1621) <= '1' when (V_X_CTRL_ANNUL_shadow /= R.X.CTRL.ANNUL) else '0';
dfp_trap_vector(1622) <= '1' when (V_X_CTRL_ANNUL_shadow /= R_A_CTRL_ANNUL_intermed_2) else '0';
dfp_trap_vector(1623) <= '1' when (V_X_CTRL_ANNUL_shadow /= V_M_CTRL_ANNUL_shadow_intermed_1) else '0';
dfp_trap_vector(1624) <= '1' when (V_X_CTRL_ANNUL_shadow /= R_X_ANNUL_ALL_intermed_1) else '0';
dfp_trap_vector(1625) <= '1' when (V_X_CTRL_ANNUL_shadow /= R.M.CTRL.ANNUL) else '0';
dfp_trap_vector(1626) <= '1' when (V_X_CTRL_ANNUL_shadow /= RIN_X_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(1627) <= '1' when (V_X_CTRL_ANNUL_shadow /= '1') else '0';
dfp_trap_vector(1628) <= '1' when (V_X_CTRL_ANNUL_shadow /= '0') else '0';
dfp_trap_vector(1629) <= '1' when (V_X_CTRL_ANNUL_shadow /= RIN_M_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(1630) <= '1' when (V_X_CTRL_ANNUL_shadow /= V_X_ANNUL_ALL_shadow_intermed_1) else '0';
dfp_trap_vector(1631) <= '1' when (V_X_CTRL_ANNUL_shadow /= RIN_E_CTRL_ANNUL_intermed_2) else '0';
dfp_trap_vector(1632) <= '1' when (V_X_CTRL_ANNUL_shadow /= RIN_X_ANNUL_ALL_intermed_2) else '0';
dfp_trap_vector(1633) <= '1' when (V_X_CTRL_ANNUL_shadow /= V_E_CTRL_ANNUL_shadow_intermed_2) else '0';
dfp_trap_vector(1634) <= '1' when (V_X_CTRL_ANNUL_shadow /= V_A_CTRL_ANNUL_shadow_intermed_3) else '0';
dfp_trap_vector(1635) <= '1' when (V_X_CTRL_ANNUL_shadow /= R_E_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(1636) <= '1' when (V_X_CTRL_TT_shadow /= V_E_CTRL_TT_shadow_intermed_3) else '0';
dfp_trap_vector(1637) <= '1' when (V_X_CTRL_TT_shadow /= RIN_A_CTRL_TT_intermed_4) else '0';
dfp_trap_vector(1638) <= '1' when (V_X_CTRL_TT_shadow /= R_A_CTRL_TT_intermed_3) else '0';
dfp_trap_vector(1639) <= '1' when (V_X_CTRL_TT_shadow /= R_M_CTRL_TT_intermed_1) else '0';
dfp_trap_vector(1640) <= '1' when (V_X_CTRL_TT_shadow /= "000000") else '0';
dfp_trap_vector(1641) <= '1' when (V_X_CTRL_TT_shadow /= R_E_CTRL_TT_intermed_2) else '0';
dfp_trap_vector(1642) <= '1' when (V_X_CTRL_TT_shadow /= R.X.CTRL.TT) else '0';
dfp_trap_vector(1643) <= '1' when (V_X_CTRL_TT_shadow /= RIN_M_CTRL_TT_intermed_2) else '0';
dfp_trap_vector(1644) <= '1' when (V_X_CTRL_TT_shadow /= RIN_E_CTRL_TT_intermed_3) else '0';
dfp_trap_vector(1645) <= '1' when (V_X_CTRL_TT_shadow /= V_M_CTRL_TT_shadow_intermed_2) else '0';
dfp_trap_vector(1646) <= '1' when (V_X_CTRL_TT_shadow /= V_A_CTRL_TT_shadow_intermed_4) else '0';
dfp_trap_vector(1647) <= '1' when (V_X_CTRL_TT_shadow /= RIN_X_CTRL_TT_intermed_1) else '0';
dfp_trap_vector(1648) <= '1' when (V_X_DATA0_shadow /= R.X.DATA ( 0 )) else '0';
dfp_trap_vector(1649) <= '1' when (V_X_DATA0_shadow /= DCO.DATA ( 0 )) else '0';
dfp_trap_vector(1650) <= '1' when (V_X_DATA0_shadow /= V_X_DATA0_shadow_intermed_2) else '0';
dfp_trap_vector(1651) <= '1' when (V_X_DATA0_shadow /= RIN_X_DATA0_intermed_1) else '0';
dfp_trap_vector(1652) <= '1' when (V_X_DATA0_shadow /= R_X_DATA0_intermed_1) else '0';
dfp_trap_vector(1653) <= '1' when (V_X_DATA0_shadow /= RIN_X_DATA0_intermed_2) else '0';
dfp_trap_vector(1654) <= '1' when (V_X_DATA1_shadow /= DCO.DATA ( 1 )) else '0';
dfp_trap_vector(1655) <= '1' when (V_X_DATA1_shadow /= R.X.DATA ( 1 )) else '0';
dfp_trap_vector(1656) <= '1' when (V_X_DATA1_shadow /= V_X_DATA1_shadow_intermed_2) else '0';
dfp_trap_vector(1657) <= '1' when (V_X_DATA1_shadow /= RIN_X_DATA1_intermed_1) else '0';
dfp_trap_vector(1658) <= '1' when (V_X_DATA1_shadow /= R_X_DATA1_intermed_1) else '0';
dfp_trap_vector(1659) <= '1' when (V_X_DATA1_shadow /= RIN_X_DATA1_intermed_2) else '0';
dfp_trap_vector(1660) <= '1' when (V_X_SET_shadow /= RIN_X_SET_intermed_1) else '0';
dfp_trap_vector(1661) <= '1' when (V_X_SET_shadow /= DCO.SET ( 0 DOWNTO 0 )) else '0';
dfp_trap_vector(1662) <= '1' when (V_X_SET_shadow /= R.X.SET) else '0';
dfp_trap_vector(1663) <= '1' when (V_X_DCI_SIZE_shadow /= R.X.DCI.SIZE) else '0';
dfp_trap_vector(1664) <= '1' when (V_X_DCI_SIZE_shadow /= V_M_DCI_SIZE_shadow_intermed_2) else '0';
dfp_trap_vector(1665) <= '1' when (V_X_DCI_SIZE_shadow /= R_M_DCI_SIZE_intermed_1) else '0';
dfp_trap_vector(1666) <= '1' when (V_X_DCI_SIZE_shadow /= RIN_X_DCI_SIZE_intermed_1) else '0';
dfp_trap_vector(1667) <= '1' when (V_X_DCI_SIZE_shadow /= RIN_M_DCI_SIZE_intermed_2) else '0';
dfp_trap_vector(1668) <= '1' when (V_X_DCI_SIGNED_shadow /= RIN_M_DCI_SIGNED_intermed_2) else '0';
dfp_trap_vector(1669) <= '1' when (V_X_DCI_SIGNED_shadow /= R_M_DCI_SIGNED_intermed_1) else '0';
dfp_trap_vector(1670) <= '1' when (V_X_DCI_SIGNED_shadow /= RIN_X_DCI_SIGNED_intermed_1) else '0';
dfp_trap_vector(1671) <= '1' when (V_X_DCI_SIGNED_shadow /= V_M_DCI_SIGNED_shadow_intermed_2) else '0';
dfp_trap_vector(1672) <= '1' when (V_X_DCI_SIGNED_shadow /= R.X.DCI.SIGNED) else '0';
dfp_trap_vector(1673) <= '1' when (V_X_MEXC_shadow /= R.X.MEXC) else '0';
dfp_trap_vector(1674) <= '1' when (V_X_MEXC_shadow /= RIN_X_MEXC_intermed_1) else '0';
dfp_trap_vector(1675) <= '1' when (V_X_MEXC_shadow /= DCO.MEXC) else '0';
dfp_trap_vector(1676) <= '1' when (V_X_ICC_shadow /= R.X.ICC) else '0';
dfp_trap_vector(1677) <= '1' when (V_X_ICC_shadow /= RIN_X_ICC_intermed_1) else '0';
dfp_trap_vector(1678) <= '1' when (V_X_ICC_shadow /= ME_ICC_shadow) else '0';
dfp_trap_vector(1679) <= '1' when (V_X_CTRL_WICC_shadow /= R_A_CTRL_WICC_intermed_2) else '0';
dfp_trap_vector(1680) <= '1' when (V_X_CTRL_WICC_shadow /= RIN_A_CTRL_ANNUL_intermed_4) else '0';
dfp_trap_vector(1681) <= '1' when (V_X_CTRL_WICC_shadow /= V_E_CTRL_WICC_shadow_intermed_2) else '0';
dfp_trap_vector(1682) <= '1' when (V_X_CTRL_WICC_shadow /= R.M.CTRL.WICC) else '0';
dfp_trap_vector(1683) <= '1' when (V_X_CTRL_WICC_shadow /= V_A_CTRL_WICC_shadow_intermed_3) else '0';
dfp_trap_vector(1684) <= '1' when (V_X_CTRL_WICC_shadow /= R_A_CTRL_ANNUL_intermed_3) else '0';
dfp_trap_vector(1685) <= '1' when (V_X_CTRL_WICC_shadow /= RIN_X_CTRL_WICC_intermed_1) else '0';
dfp_trap_vector(1686) <= '1' when (V_X_CTRL_WICC_shadow /= R_X_ANNUL_ALL_intermed_3) else '0';
dfp_trap_vector(1687) <= '1' when (V_X_CTRL_WICC_shadow /= RIN_E_CTRL_WICC_intermed_2) else '0';
dfp_trap_vector(1688) <= '1' when (V_X_CTRL_WICC_shadow /= RIN_M_CTRL_WICC_intermed_1) else '0';
dfp_trap_vector(1689) <= '1' when (V_X_CTRL_WICC_shadow /= R.X.CTRL.WICC) else '0';
dfp_trap_vector(1690) <= '1' when (V_X_CTRL_WICC_shadow /= '1') else '0';
dfp_trap_vector(1691) <= '1' when (V_X_CTRL_WICC_shadow /= '0') else '0';
dfp_trap_vector(1692) <= '1' when (V_X_CTRL_WICC_shadow /= R_E_CTRL_WICC_intermed_1) else '0';
dfp_trap_vector(1693) <= '1' when (V_X_CTRL_WICC_shadow /= V_X_ANNUL_ALL_shadow_intermed_3) else '0';
dfp_trap_vector(1694) <= '1' when (V_X_CTRL_WICC_shadow /= V_M_CTRL_WICC_shadow_intermed_1) else '0';
dfp_trap_vector(1695) <= '1' when (V_X_CTRL_WICC_shadow /= RIN_X_ANNUL_ALL_intermed_4) else '0';
dfp_trap_vector(1696) <= '1' when (V_X_CTRL_WICC_shadow /= RIN_A_CTRL_WICC_intermed_3) else '0';
dfp_trap_vector(1697) <= '1' when (V_X_CTRL_WICC_shadow /= V_A_CTRL_ANNUL_shadow_intermed_3) else '0';
dfp_trap_vector(1698) <= '1' when (V_M_CTRL_shadow /= RIN_E_CTRL_intermed_1) else '0';
dfp_trap_vector(1699) <= '1' when (V_M_CTRL_shadow /= R.E.CTRL) else '0';
dfp_trap_vector(1700) <= '1' when (V_M_CTRL_shadow /= R.M.CTRL) else '0';
dfp_trap_vector(1701) <= '1' when (V_M_CTRL_shadow /= RIN_M_CTRL_intermed_1) else '0';
dfp_trap_vector(1702) <= '1' when (V_M_CTRL_shadow /= V_E_CTRL_shadow_intermed_1) else '0';
dfp_trap_vector(1703) <= '1' when (V_M_CTRL_shadow /= RIN_A_CTRL_intermed_2) else '0';
dfp_trap_vector(1704) <= '1' when (V_M_CTRL_shadow /= V_A_CTRL_shadow_intermed_2) else '0';
dfp_trap_vector(1705) <= '1' when (V_M_CTRL_shadow /= R_A_CTRL_intermed_1) else '0';
dfp_trap_vector(1706) <= '1' when (V_M_CTRL_RETT_shadow /= R.M.CTRL.RETT) else '0';
dfp_trap_vector(1707) <= '1' when (V_M_CTRL_RETT_shadow /= RIN_A_CTRL_ANNUL_intermed_3) else '0';
dfp_trap_vector(1708) <= '1' when (V_M_CTRL_RETT_shadow /= R_A_CTRL_ANNUL_intermed_2) else '0';
dfp_trap_vector(1709) <= '1' when (V_M_CTRL_RETT_shadow /= RIN_M_CTRL_RETT_intermed_1) else '0';
dfp_trap_vector(1710) <= '1' when (V_M_CTRL_RETT_shadow /= R_X_ANNUL_ALL_intermed_2) else '0';
dfp_trap_vector(1711) <= '1' when (V_M_CTRL_RETT_shadow /= '1') else '0';
dfp_trap_vector(1712) <= '1' when (V_M_CTRL_RETT_shadow /= '0') else '0';
dfp_trap_vector(1713) <= '1' when (V_M_CTRL_RETT_shadow /= V_E_CTRL_RETT_shadow_intermed_1) else '0';
dfp_trap_vector(1714) <= '1' when (V_M_CTRL_RETT_shadow /= V_A_CTRL_RETT_shadow_intermed_2) else '0';
dfp_trap_vector(1715) <= '1' when (V_M_CTRL_RETT_shadow /= RIN_A_CTRL_RETT_intermed_2) else '0';
dfp_trap_vector(1716) <= '1' when (V_M_CTRL_RETT_shadow /= V_X_ANNUL_ALL_shadow_intermed_2) else '0';
dfp_trap_vector(1717) <= '1' when (V_M_CTRL_RETT_shadow /= RIN_E_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(1718) <= '1' when (V_M_CTRL_RETT_shadow /= R.E.CTRL.RETT) else '0';
dfp_trap_vector(1719) <= '1' when (V_M_CTRL_RETT_shadow /= RIN_X_ANNUL_ALL_intermed_3) else '0';
dfp_trap_vector(1720) <= '1' when (V_M_CTRL_RETT_shadow /= RIN_E_CTRL_RETT_intermed_1) else '0';
dfp_trap_vector(1721) <= '1' when (V_M_CTRL_RETT_shadow /= V_E_CTRL_ANNUL_shadow_intermed_1) else '0';
dfp_trap_vector(1722) <= '1' when (V_M_CTRL_RETT_shadow /= V_A_CTRL_ANNUL_shadow_intermed_2) else '0';
dfp_trap_vector(1723) <= '1' when (V_M_CTRL_RETT_shadow /= R_A_CTRL_RETT_intermed_1) else '0';
dfp_trap_vector(1724) <= '1' when (V_M_CTRL_RETT_shadow /= R.E.CTRL.ANNUL) else '0';
dfp_trap_vector(1725) <= '1' when (V_M_CTRL_WREG_shadow /= RIN_A_CTRL_ANNUL_intermed_3) else '0';
dfp_trap_vector(1726) <= '1' when (V_M_CTRL_WREG_shadow /= R_A_CTRL_ANNUL_intermed_2) else '0';
dfp_trap_vector(1727) <= '1' when (V_M_CTRL_WREG_shadow /= R_X_ANNUL_ALL_intermed_2) else '0';
dfp_trap_vector(1728) <= '1' when (V_M_CTRL_WREG_shadow /= '1') else '0';
dfp_trap_vector(1729) <= '1' when (V_M_CTRL_WREG_shadow /= '0') else '0';
dfp_trap_vector(1730) <= '1' when (V_M_CTRL_WREG_shadow /= RIN_M_CTRL_WREG_intermed_1) else '0';
dfp_trap_vector(1731) <= '1' when (V_M_CTRL_WREG_shadow /= RIN_A_CTRL_WREG_intermed_2) else '0';
dfp_trap_vector(1732) <= '1' when (V_M_CTRL_WREG_shadow /= V_A_CTRL_WREG_shadow_intermed_2) else '0';
dfp_trap_vector(1733) <= '1' when (V_M_CTRL_WREG_shadow /= R_A_CTRL_WREG_intermed_1) else '0';
dfp_trap_vector(1734) <= '1' when (V_M_CTRL_WREG_shadow /= V_X_ANNUL_ALL_shadow_intermed_2) else '0';
dfp_trap_vector(1735) <= '1' when (V_M_CTRL_WREG_shadow /= R.M.CTRL.WREG) else '0';
dfp_trap_vector(1736) <= '1' when (V_M_CTRL_WREG_shadow /= RIN_X_ANNUL_ALL_intermed_3) else '0';
dfp_trap_vector(1737) <= '1' when (V_M_CTRL_WREG_shadow /= R.E.CTRL.WREG) else '0';
dfp_trap_vector(1738) <= '1' when (V_M_CTRL_WREG_shadow /= V_A_CTRL_ANNUL_shadow_intermed_2) else '0';
dfp_trap_vector(1739) <= '1' when (V_M_CTRL_WREG_shadow /= RIN_E_CTRL_WREG_intermed_1) else '0';
dfp_trap_vector(1740) <= '1' when (V_M_CTRL_WREG_shadow /= V_E_CTRL_WREG_shadow_intermed_1) else '0';
dfp_trap_vector(1741) <= '1' when (V_E_CWP_shadow /= RIN_E_CWP_intermed_1) else '0';
dfp_trap_vector(1742) <= '1' when (V_E_CWP_shadow /= V_A_CWP_shadow_intermed_1) else '0';
dfp_trap_vector(1743) <= '1' when (V_E_CWP_shadow /= RIN_D_CWP_intermed_2) else '0';
dfp_trap_vector(1744) <= '1' when (V_E_CWP_shadow /= R.E.CWP) else '0';
dfp_trap_vector(1745) <= '1' when (V_E_CWP_shadow /= RIN_A_CWP_intermed_1) else '0';
dfp_trap_vector(1746) <= '1' when (V_E_CWP_shadow /= V_D_CWP_shadow_intermed_2) else '0';
dfp_trap_vector(1747) <= '1' when (V_E_CWP_shadow /= R_D_CWP_intermed_1) else '0';
dfp_trap_vector(1748) <= '1' when (V_E_CWP_shadow /= R.A.CWP) else '0';
dfp_trap_vector(1749) <= '1' when (V_M_SU_shadow /= R.M.SU) else '0';
dfp_trap_vector(1750) <= '1' when (V_M_SU_shadow /= R_A_SU_intermed_1) else '0';
dfp_trap_vector(1751) <= '1' when (V_M_SU_shadow /= RIN_A_SU_intermed_2) else '0';
dfp_trap_vector(1752) <= '1' when (V_M_SU_shadow /= V_E_SU_shadow_intermed_1) else '0';
dfp_trap_vector(1753) <= '1' when (V_M_SU_shadow /= R.E.SU) else '0';
dfp_trap_vector(1754) <= '1' when (V_M_SU_shadow /= V_A_SU_shadow_intermed_2) else '0';
dfp_trap_vector(1755) <= '1' when (V_M_SU_shadow /= RIN_M_SU_intermed_1) else '0';
dfp_trap_vector(1756) <= '1' when (V_M_SU_shadow /= RIN_E_SU_intermed_1) else '0';
dfp_trap_vector(1757) <= '1' when (V_M_MUL_shadow /= RIN_M_MUL_intermed_1) else '0';
dfp_trap_vector(1758) <= '1' when (V_M_MUL_shadow /= '0') else '0';
dfp_trap_vector(1759) <= '1' when (V_M_MUL_shadow /= R.M.MUL) else '0';
dfp_trap_vector(1760) <= '1' when (V_M_NALIGN_shadow /= '1') else '0';
dfp_trap_vector(1761) <= '1' when (V_M_NALIGN_shadow /= '0') else '0';
dfp_trap_vector(1762) <= '1' when (V_M_NALIGN_shadow /= RIN_M_NALIGN_intermed_1) else '0';
dfp_trap_vector(1763) <= '1' when (V_M_NALIGN_shadow /= R.M.NALIGN) else '0';
dfp_trap_vector(1764) <= '1' when (EX_ADD_RES3_shadow /= EX_OP23_shadow) else '0';
dfp_trap_vector(1765) <= '1' when (EX_ADD_RES3_shadow /= V_X_DATA03_shadow_intermed_2) else '0';
dfp_trap_vector(1766) <= '1' when (EX_ADD_RES3_shadow /= V_X_DATA03_shadow_intermed_1) else '0';
dfp_trap_vector(1767) <= '1' when (EX_ADD_RES3_shadow /= DCO_DATA03_intermed_1) else '0';
dfp_trap_vector(1768) <= '1' when (EX_ADD_RES3_shadow /= R.E.OP2( 3 )) else '0';
dfp_trap_vector(1769) <= '1' when (EX_ADD_RES3_shadow /= RIN_X_DATA03_intermed_1) else '0';
dfp_trap_vector(1770) <= '1' when (EX_ADD_RES3_shadow /= R_X_DATA03_intermed_1) else '0';
dfp_trap_vector(1771) <= '1' when (EX_ADD_RES3_shadow /= RIN_X_DATA03_intermed_2) else '0';
dfp_trap_vector(1772) <= '1' when (EX_ADD_RES3_shadow /= RIN_E_OP23_intermed_1) else '0';
dfp_trap_vector(1773) <= '1' when (EX_ADD_RES3_shadow /= RIN_E_OP13_intermed_1) else '0';
dfp_trap_vector(1774) <= '1' when (EX_ADD_RES3_shadow /= EX_FORCE_A2_shadow) else '0';
dfp_trap_vector(1775) <= '1' when (EX_ADD_RES3_shadow /= R.X.DATA ( 0 )( 3 )) else '0';
dfp_trap_vector(1776) <= '1' when (EX_ADD_RES3_shadow /= EX_OP13_shadow) else '0';
dfp_trap_vector(1777) <= '1' when (EX_ADD_RES3_shadow /= V_E_OP23_shadow_intermed_1) else '0';
dfp_trap_vector(1778) <= '1' when (EX_ADD_RES3_shadow /= R.E.OP1( 3 )) else '0';
dfp_trap_vector(1779) <= '1' when (EX_ADD_RES3_shadow /= V_E_OP13_shadow_intermed_1) else '0';
dfp_trap_vector(1780) <= '1' when (V_M_CTRL_ANNUL_shadow /= RIN_A_CTRL_ANNUL_intermed_3) else '0';
dfp_trap_vector(1781) <= '1' when (V_M_CTRL_ANNUL_shadow /= R_A_CTRL_ANNUL_intermed_2) else '0';
dfp_trap_vector(1782) <= '1' when (V_M_CTRL_ANNUL_shadow /= R.X.ANNUL_ALL) else '0';
dfp_trap_vector(1783) <= '1' when (V_M_CTRL_ANNUL_shadow /= R.M.CTRL.ANNUL) else '0';
dfp_trap_vector(1784) <= '1' when (V_M_CTRL_ANNUL_shadow /= '1') else '0';
dfp_trap_vector(1785) <= '1' when (V_M_CTRL_ANNUL_shadow /= '0') else '0';
dfp_trap_vector(1786) <= '1' when (V_M_CTRL_ANNUL_shadow /= RIN_M_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(1787) <= '1' when (V_M_CTRL_ANNUL_shadow /= V_X_ANNUL_ALL_shadow) else '0';
dfp_trap_vector(1788) <= '1' when (V_M_CTRL_ANNUL_shadow /= RIN_E_CTRL_ANNUL_intermed_2) else '0';
dfp_trap_vector(1789) <= '1' when (V_M_CTRL_ANNUL_shadow /= RIN_X_ANNUL_ALL_intermed_1) else '0';
dfp_trap_vector(1790) <= '1' when (V_M_CTRL_ANNUL_shadow /= V_E_CTRL_ANNUL_shadow_intermed_2) else '0';
dfp_trap_vector(1791) <= '1' when (V_M_CTRL_ANNUL_shadow /= V_A_CTRL_ANNUL_shadow_intermed_3) else '0';
dfp_trap_vector(1792) <= '1' when (V_M_CTRL_ANNUL_shadow /= R_E_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(1793) <= '1' when (V_M_CTRL_WICC_shadow /= R_A_CTRL_WICC_intermed_1) else '0';
dfp_trap_vector(1794) <= '1' when (V_M_CTRL_WICC_shadow /= RIN_A_CTRL_ANNUL_intermed_3) else '0';
dfp_trap_vector(1795) <= '1' when (V_M_CTRL_WICC_shadow /= V_E_CTRL_WICC_shadow_intermed_1) else '0';
dfp_trap_vector(1796) <= '1' when (V_M_CTRL_WICC_shadow /= R.M.CTRL.WICC) else '0';
dfp_trap_vector(1797) <= '1' when (V_M_CTRL_WICC_shadow /= V_A_CTRL_WICC_shadow_intermed_2) else '0';
dfp_trap_vector(1798) <= '1' when (V_M_CTRL_WICC_shadow /= R_A_CTRL_ANNUL_intermed_2) else '0';
dfp_trap_vector(1799) <= '1' when (V_M_CTRL_WICC_shadow /= R_X_ANNUL_ALL_intermed_2) else '0';
dfp_trap_vector(1800) <= '1' when (V_M_CTRL_WICC_shadow /= RIN_E_CTRL_WICC_intermed_1) else '0';
dfp_trap_vector(1801) <= '1' when (V_M_CTRL_WICC_shadow /= RIN_M_CTRL_WICC_intermed_1) else '0';
dfp_trap_vector(1802) <= '1' when (V_M_CTRL_WICC_shadow /= '1') else '0';
dfp_trap_vector(1803) <= '1' when (V_M_CTRL_WICC_shadow /= '0') else '0';
dfp_trap_vector(1804) <= '1' when (V_M_CTRL_WICC_shadow /= R.E.CTRL.WICC) else '0';
dfp_trap_vector(1805) <= '1' when (V_M_CTRL_WICC_shadow /= V_X_ANNUL_ALL_shadow_intermed_2) else '0';
dfp_trap_vector(1806) <= '1' when (V_M_CTRL_WICC_shadow /= RIN_X_ANNUL_ALL_intermed_3) else '0';
dfp_trap_vector(1807) <= '1' when (V_M_CTRL_WICC_shadow /= RIN_A_CTRL_WICC_intermed_2) else '0';
dfp_trap_vector(1808) <= '1' when (V_M_CTRL_WICC_shadow /= V_A_CTRL_ANNUL_shadow_intermed_2) else '0';
dfp_trap_vector(1809) <= '1' when (V_M_MAC_shadow /= V_E_MAC_shadow_intermed_1) else '0';
dfp_trap_vector(1810) <= '1' when (V_M_MAC_shadow /= RIN_M_MAC_intermed_1) else '0';
dfp_trap_vector(1811) <= '1' when (V_M_MAC_shadow /= RIN_E_MAC_intermed_1) else '0';
dfp_trap_vector(1812) <= '1' when (V_M_MAC_shadow /= R.E.MAC) else '0';
dfp_trap_vector(1813) <= '1' when (V_M_MAC_shadow /= R.M.MAC) else '0';
dfp_trap_vector(1814) <= '1' when (V_M_CTRL_LD_shadow /= R_A_CTRL_LD_intermed_2) else '0';
dfp_trap_vector(1815) <= '1' when (V_M_CTRL_LD_shadow /= RIN_A_CTRL_LD_intermed_3) else '0';
dfp_trap_vector(1816) <= '1' when (V_M_CTRL_LD_shadow /= V_E_CTRL_LD_shadow_intermed_2) else '0';
dfp_trap_vector(1817) <= '1' when (V_M_CTRL_LD_shadow /= '1') else '0';
dfp_trap_vector(1818) <= '1' when (V_M_CTRL_LD_shadow /= R_E_CTRL_LD_intermed_1) else '0';
dfp_trap_vector(1819) <= '1' when (V_M_CTRL_LD_shadow /= R.M.CTRL.LD) else '0';
dfp_trap_vector(1820) <= '1' when (V_M_CTRL_LD_shadow /= RIN_E_CTRL_LD_intermed_2) else '0';
dfp_trap_vector(1821) <= '1' when (V_M_CTRL_LD_shadow /= RIN_M_CTRL_LD_intermed_1) else '0';
dfp_trap_vector(1822) <= '1' when (V_M_CTRL_LD_shadow /= V_A_CTRL_LD_shadow_intermed_3) else '0';
dfp_trap_vector(1823) <= '1' when (V_E_CTRL_shadow /= RIN_E_CTRL_intermed_1) else '0';
dfp_trap_vector(1824) <= '1' when (V_E_CTRL_shadow /= R.E.CTRL) else '0';
dfp_trap_vector(1825) <= '1' when (V_E_CTRL_shadow /= RIN_A_CTRL_intermed_1) else '0';
dfp_trap_vector(1826) <= '1' when (V_E_CTRL_shadow /= V_A_CTRL_shadow_intermed_1) else '0';
dfp_trap_vector(1827) <= '1' when (V_E_CTRL_shadow /= R.A.CTRL) else '0';
dfp_trap_vector(1828) <= '1' when (V_E_JMPL_shadow /= RIN_E_JMPL_intermed_1) else '0';
dfp_trap_vector(1829) <= '1' when (V_E_JMPL_shadow /= R.A.JMPL) else '0';
dfp_trap_vector(1830) <= '1' when (V_E_JMPL_shadow /= RIN_A_JMPL_intermed_1) else '0';
dfp_trap_vector(1831) <= '1' when (V_E_JMPL_shadow /= R.E.JMPL) else '0';
dfp_trap_vector(1832) <= '1' when (V_E_JMPL_shadow /= V_A_JMPL_shadow_intermed_1) else '0';
dfp_trap_vector(1833) <= '1' when (V_E_CTRL_ANNUL_shadow /= RIN_A_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(1834) <= '1' when (V_E_CTRL_ANNUL_shadow /= R.A.CTRL.ANNUL) else '0';
dfp_trap_vector(1835) <= '1' when (V_E_CTRL_ANNUL_shadow /= R_X_ANNUL_ALL_intermed_1) else '0';
dfp_trap_vector(1836) <= '1' when (V_E_CTRL_ANNUL_shadow /= '1') else '0';
dfp_trap_vector(1837) <= '1' when (V_E_CTRL_ANNUL_shadow /= '0') else '0';
dfp_trap_vector(1838) <= '1' when (V_E_CTRL_ANNUL_shadow /= V_X_ANNUL_ALL_shadow_intermed_1) else '0';
dfp_trap_vector(1839) <= '1' when (V_E_CTRL_ANNUL_shadow /= RIN_E_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(1840) <= '1' when (V_E_CTRL_ANNUL_shadow /= RIN_X_ANNUL_ALL_intermed_2) else '0';
dfp_trap_vector(1841) <= '1' when (V_E_CTRL_ANNUL_shadow /= V_A_CTRL_ANNUL_shadow_intermed_1) else '0';
dfp_trap_vector(1842) <= '1' when (V_E_CTRL_ANNUL_shadow /= R.E.CTRL.ANNUL) else '0';
dfp_trap_vector(1843) <= '1' when (V_E_CTRL_RETT_shadow /= RIN_A_CTRL_ANNUL_intermed_2) else '0';
dfp_trap_vector(1844) <= '1' when (V_E_CTRL_RETT_shadow /= R_A_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(1845) <= '1' when (V_E_CTRL_RETT_shadow /= R_X_ANNUL_ALL_intermed_1) else '0';
dfp_trap_vector(1846) <= '1' when (V_E_CTRL_RETT_shadow /= '1') else '0';
dfp_trap_vector(1847) <= '1' when (V_E_CTRL_RETT_shadow /= '0') else '0';
dfp_trap_vector(1848) <= '1' when (V_E_CTRL_RETT_shadow /= V_A_CTRL_RETT_shadow_intermed_1) else '0';
dfp_trap_vector(1849) <= '1' when (V_E_CTRL_RETT_shadow /= RIN_A_CTRL_RETT_intermed_1) else '0';
dfp_trap_vector(1850) <= '1' when (V_E_CTRL_RETT_shadow /= V_X_ANNUL_ALL_shadow_intermed_1) else '0';
dfp_trap_vector(1851) <= '1' when (V_E_CTRL_RETT_shadow /= R.E.CTRL.RETT) else '0';
dfp_trap_vector(1852) <= '1' when (V_E_CTRL_RETT_shadow /= RIN_X_ANNUL_ALL_intermed_2) else '0';
dfp_trap_vector(1853) <= '1' when (V_E_CTRL_RETT_shadow /= RIN_E_CTRL_RETT_intermed_1) else '0';
dfp_trap_vector(1854) <= '1' when (V_E_CTRL_RETT_shadow /= V_A_CTRL_ANNUL_shadow_intermed_1) else '0';
dfp_trap_vector(1855) <= '1' when (V_E_CTRL_RETT_shadow /= R.A.CTRL.RETT) else '0';
dfp_trap_vector(1856) <= '1' when (V_E_CTRL_WREG_shadow /= RIN_A_CTRL_ANNUL_intermed_2) else '0';
dfp_trap_vector(1857) <= '1' when (V_E_CTRL_WREG_shadow /= R_A_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(1858) <= '1' when (V_E_CTRL_WREG_shadow /= R_X_ANNUL_ALL_intermed_1) else '0';
dfp_trap_vector(1859) <= '1' when (V_E_CTRL_WREG_shadow /= '1') else '0';
dfp_trap_vector(1860) <= '1' when (V_E_CTRL_WREG_shadow /= '0') else '0';
dfp_trap_vector(1861) <= '1' when (V_E_CTRL_WREG_shadow /= RIN_A_CTRL_WREG_intermed_1) else '0';
dfp_trap_vector(1862) <= '1' when (V_E_CTRL_WREG_shadow /= V_A_CTRL_WREG_shadow_intermed_1) else '0';
dfp_trap_vector(1863) <= '1' when (V_E_CTRL_WREG_shadow /= R.A.CTRL.WREG) else '0';
dfp_trap_vector(1864) <= '1' when (V_E_CTRL_WREG_shadow /= V_X_ANNUL_ALL_shadow_intermed_1) else '0';
dfp_trap_vector(1865) <= '1' when (V_E_CTRL_WREG_shadow /= RIN_X_ANNUL_ALL_intermed_2) else '0';
dfp_trap_vector(1866) <= '1' when (V_E_CTRL_WREG_shadow /= R.E.CTRL.WREG) else '0';
dfp_trap_vector(1867) <= '1' when (V_E_CTRL_WREG_shadow /= V_A_CTRL_ANNUL_shadow_intermed_1) else '0';
dfp_trap_vector(1868) <= '1' when (V_E_CTRL_WREG_shadow /= RIN_E_CTRL_WREG_intermed_1) else '0';
dfp_trap_vector(1869) <= '1' when (V_E_SU_shadow /= R.A.SU) else '0';
dfp_trap_vector(1870) <= '1' when (V_E_SU_shadow /= RIN_A_SU_intermed_1) else '0';
dfp_trap_vector(1871) <= '1' when (V_E_SU_shadow /= R.E.SU) else '0';
dfp_trap_vector(1872) <= '1' when (V_E_SU_shadow /= V_A_SU_shadow_intermed_1) else '0';
dfp_trap_vector(1873) <= '1' when (V_E_SU_shadow /= RIN_E_SU_intermed_1) else '0';
dfp_trap_vector(1874) <= '1' when (V_E_ET_shadow /= RIN_E_ET_intermed_1) else '0';
dfp_trap_vector(1875) <= '1' when (V_E_ET_shadow /= R.E.ET) else '0';
dfp_trap_vector(1876) <= '1' when (V_E_ET_shadow /= RIN_A_ET_intermed_1) else '0';
dfp_trap_vector(1877) <= '1' when (V_E_ET_shadow /= V_A_ET_shadow_intermed_1) else '0';
dfp_trap_vector(1878) <= '1' when (V_E_ET_shadow /= R.A.ET) else '0';
dfp_trap_vector(1879) <= '1' when (V_E_CTRL_WICC_shadow /= R.A.CTRL.WICC) else '0';
dfp_trap_vector(1880) <= '1' when (V_E_CTRL_WICC_shadow /= RIN_A_CTRL_ANNUL_intermed_2) else '0';
dfp_trap_vector(1881) <= '1' when (V_E_CTRL_WICC_shadow /= V_A_CTRL_WICC_shadow_intermed_1) else '0';
dfp_trap_vector(1882) <= '1' when (V_E_CTRL_WICC_shadow /= R_A_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(1883) <= '1' when (V_E_CTRL_WICC_shadow /= RIN_E_CTRL_WICC_intermed_1) else '0';
dfp_trap_vector(1884) <= '1' when (V_E_CTRL_WICC_shadow /= R_X_ANNUL_ALL_intermed_1) else '0';
dfp_trap_vector(1885) <= '1' when (V_E_CTRL_WICC_shadow /= '1') else '0';
dfp_trap_vector(1886) <= '1' when (V_E_CTRL_WICC_shadow /= '0') else '0';
dfp_trap_vector(1887) <= '1' when (V_E_CTRL_WICC_shadow /= R.E.CTRL.WICC) else '0';
dfp_trap_vector(1888) <= '1' when (V_E_CTRL_WICC_shadow /= V_X_ANNUL_ALL_shadow_intermed_1) else '0';
dfp_trap_vector(1889) <= '1' when (V_E_CTRL_WICC_shadow /= RIN_X_ANNUL_ALL_intermed_2) else '0';
dfp_trap_vector(1890) <= '1' when (V_E_CTRL_WICC_shadow /= RIN_A_CTRL_WICC_intermed_1) else '0';
dfp_trap_vector(1891) <= '1' when (V_E_CTRL_WICC_shadow /= V_A_CTRL_ANNUL_shadow_intermed_1) else '0';
dfp_trap_vector(1892) <= '1' when (V_A_CWP_shadow /= RIN_D_CWP_intermed_1) else '0';
dfp_trap_vector(1893) <= '1' when (V_A_CWP_shadow /= RIN_A_CWP_intermed_1) else '0';
dfp_trap_vector(1894) <= '1' when (V_A_CWP_shadow /= V_D_CWP_shadow_intermed_1) else '0';
dfp_trap_vector(1895) <= '1' when (V_A_CWP_shadow /= R.D.CWP) else '0';
dfp_trap_vector(1896) <= '1' when (V_A_CWP_shadow /= R.A.CWP) else '0';
dfp_trap_vector(1897) <= '1' when (V_A_RFA1_shadow /= DBGI.DADDR ( 9 DOWNTO 2 )) else '0';
dfp_trap_vector(1898) <= '1' when (V_A_RFA1_shadow /= DE_RADDR17DOWNTO0_shadow) else '0';
dfp_trap_vector(1899) <= '1' when (V_A_RFA1_shadow /= R.A.RFA1) else '0';
dfp_trap_vector(1900) <= '1' when (V_A_RFA1_shadow /= RIN_A_RFA1_intermed_1) else '0';
dfp_trap_vector(1901) <= '1' when (DE_RADDR17DOWNTO0_shadow /= V_A_RFA1_shadow_intermed_1) else '0';
dfp_trap_vector(1902) <= '1' when (DE_RADDR17DOWNTO0_shadow /= DBGI_DADDR9DOWNTO2_intermed_1) else '0';
dfp_trap_vector(1903) <= '1' when (DE_RADDR17DOWNTO0_shadow /= R.A.RFA1) else '0';
dfp_trap_vector(1904) <= '1' when (DE_RADDR17DOWNTO0_shadow /= RIN_A_RFA1_intermed_1) else '0';
dfp_trap_vector(1905) <= '1' when (V_A_RFA2_shadow /= DE_RADDR27DOWNTO0_shadow) else '0';
dfp_trap_vector(1906) <= '1' when (V_A_RFA2_shadow /= R.A.RFA2) else '0';
dfp_trap_vector(1907) <= '1' when (V_A_RFA2_shadow /= RIN_A_RFA2_intermed_1) else '0';
dfp_trap_vector(1908) <= '1' when (V_A_CTRL_ANNUL_shadow /= RIN_A_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(1909) <= '1' when (V_A_CTRL_ANNUL_shadow /= R.A.CTRL.ANNUL) else '0';
dfp_trap_vector(1910) <= '1' when (V_A_CTRL_ANNUL_shadow /= R.X.ANNUL_ALL) else '0';
dfp_trap_vector(1911) <= '1' when (V_A_CTRL_ANNUL_shadow /= '1') else '0';
dfp_trap_vector(1912) <= '1' when (V_A_CTRL_ANNUL_shadow /= '0') else '0';
dfp_trap_vector(1913) <= '1' when (V_A_CTRL_ANNUL_shadow /= V_X_ANNUL_ALL_shadow) else '0';
dfp_trap_vector(1914) <= '1' when (V_A_CTRL_ANNUL_shadow /= RIN_X_ANNUL_ALL_intermed_1) else '0';
dfp_trap_vector(1915) <= '1' when (V_A_CTRL_WICC_shadow /= R.A.CTRL.WICC) else '0';
dfp_trap_vector(1916) <= '1' when (V_A_CTRL_WICC_shadow /= RIN_A_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(1917) <= '1' when (V_A_CTRL_WICC_shadow /= R.A.CTRL.ANNUL) else '0';
dfp_trap_vector(1918) <= '1' when (V_A_CTRL_WICC_shadow /= R.X.ANNUL_ALL) else '0';
dfp_trap_vector(1919) <= '1' when (V_A_CTRL_WICC_shadow /= '1') else '0';
dfp_trap_vector(1920) <= '1' when (V_A_CTRL_WICC_shadow /= '0') else '0';
dfp_trap_vector(1921) <= '1' when (V_A_CTRL_WICC_shadow /= V_X_ANNUL_ALL_shadow) else '0';
dfp_trap_vector(1922) <= '1' when (V_A_CTRL_WICC_shadow /= RIN_X_ANNUL_ALL_intermed_1) else '0';
dfp_trap_vector(1923) <= '1' when (V_A_CTRL_WICC_shadow /= RIN_A_CTRL_WICC_intermed_1) else '0';
dfp_trap_vector(1924) <= '1' when (V_A_CTRL_WICC_shadow /= V_A_CTRL_ANNUL_shadow) else '0';
dfp_trap_vector(1925) <= '1' when (V_A_CTRL_WREG_shadow /= RIN_A_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(1926) <= '1' when (V_A_CTRL_WREG_shadow /= R.A.CTRL.ANNUL) else '0';
dfp_trap_vector(1927) <= '1' when (V_A_CTRL_WREG_shadow /= R.X.ANNUL_ALL) else '0';
dfp_trap_vector(1928) <= '1' when (V_A_CTRL_WREG_shadow /= '1') else '0';
dfp_trap_vector(1929) <= '1' when (V_A_CTRL_WREG_shadow /= '0') else '0';
dfp_trap_vector(1930) <= '1' when (V_A_CTRL_WREG_shadow /= RIN_A_CTRL_WREG_intermed_1) else '0';
dfp_trap_vector(1931) <= '1' when (V_A_CTRL_WREG_shadow /= R.A.CTRL.WREG) else '0';
dfp_trap_vector(1932) <= '1' when (V_A_CTRL_WREG_shadow /= V_X_ANNUL_ALL_shadow) else '0';
dfp_trap_vector(1933) <= '1' when (V_A_CTRL_WREG_shadow /= RIN_X_ANNUL_ALL_intermed_1) else '0';
dfp_trap_vector(1934) <= '1' when (V_A_CTRL_WREG_shadow /= V_A_CTRL_ANNUL_shadow) else '0';
dfp_trap_vector(1935) <= '1' when (V_A_CTRL_RETT_shadow /= RIN_A_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(1936) <= '1' when (V_A_CTRL_RETT_shadow /= R.A.CTRL.ANNUL) else '0';
dfp_trap_vector(1937) <= '1' when (V_A_CTRL_RETT_shadow /= R.X.ANNUL_ALL) else '0';
dfp_trap_vector(1938) <= '1' when (V_A_CTRL_RETT_shadow /= '1') else '0';
dfp_trap_vector(1939) <= '1' when (V_A_CTRL_RETT_shadow /= '0') else '0';
dfp_trap_vector(1940) <= '1' when (V_A_CTRL_RETT_shadow /= RIN_A_CTRL_RETT_intermed_1) else '0';
dfp_trap_vector(1941) <= '1' when (V_A_CTRL_RETT_shadow /= V_X_ANNUL_ALL_shadow) else '0';
dfp_trap_vector(1942) <= '1' when (V_A_CTRL_RETT_shadow /= RIN_X_ANNUL_ALL_intermed_1) else '0';
dfp_trap_vector(1943) <= '1' when (V_A_CTRL_RETT_shadow /= V_A_CTRL_ANNUL_shadow) else '0';
dfp_trap_vector(1944) <= '1' when (V_A_CTRL_RETT_shadow /= R.A.CTRL.RETT) else '0';
dfp_trap_vector(1945) <= '1' when (V_A_CTRL_WY_shadow /= RIN_A_CTRL_ANNUL_intermed_1) else '0';
dfp_trap_vector(1946) <= '1' when (V_A_CTRL_WY_shadow /= R.A.CTRL.ANNUL) else '0';
dfp_trap_vector(1947) <= '1' when (V_A_CTRL_WY_shadow /= R.X.ANNUL_ALL) else '0';
dfp_trap_vector(1948) <= '1' when (V_A_CTRL_WY_shadow /= '1') else '0';
dfp_trap_vector(1949) <= '1' when (V_A_CTRL_WY_shadow /= '0') else '0';
dfp_trap_vector(1950) <= '1' when (V_A_CTRL_WY_shadow /= V_X_ANNUL_ALL_shadow) else '0';
dfp_trap_vector(1951) <= '1' when (V_A_CTRL_WY_shadow /= RIN_X_ANNUL_ALL_intermed_1) else '0';
dfp_trap_vector(1952) <= '1' when (V_A_CTRL_WY_shadow /= R.A.CTRL.WY) else '0';
dfp_trap_vector(1953) <= '1' when (V_A_CTRL_WY_shadow /= RIN_A_CTRL_WY_intermed_1) else '0';
dfp_trap_vector(1954) <= '1' when (V_A_CTRL_WY_shadow /= V_A_CTRL_ANNUL_shadow) else '0';
dfp_trap_vector(1955) <= '1' when (V_A_CTRL_TRAP_shadow /= ICO_MEXC_intermed_1) else '0';
dfp_trap_vector(1956) <= '1' when (V_A_CTRL_TRAP_shadow /= RIN_A_CTRL_TRAP_intermed_1) else '0';
dfp_trap_vector(1957) <= '1' when (V_A_CTRL_TRAP_shadow /= R.D.MEXC) else '0';
dfp_trap_vector(1958) <= '1' when (V_A_CTRL_TRAP_shadow /= V_D_MEXC_shadow_intermed_1) else '0';
dfp_trap_vector(1959) <= '1' when (V_A_CTRL_TRAP_shadow /= R.A.CTRL.TRAP) else '0';
dfp_trap_vector(1960) <= '1' when (V_A_CTRL_TRAP_shadow /= RIN_D_MEXC_intermed_1) else '0';
dfp_trap_vector(1961) <= '1' when (V_A_CTRL_TT_shadow /= RIN_A_CTRL_TT_intermed_1) else '0';
dfp_trap_vector(1962) <= '1' when (V_A_CTRL_TT_shadow /= R.A.CTRL.TT) else '0';
dfp_trap_vector(1963) <= '1' when (V_A_CTRL_TT_shadow /= "000000") else '0';
dfp_trap_vector(1964) <= '1' when (V_A_CTRL_INST_shadow /= DE_INST_shadow) else '0';
dfp_trap_vector(1965) <= '1' when (V_A_CTRL_INST_shadow /= RIN_A_CTRL_INST_intermed_1) else '0';
dfp_trap_vector(1966) <= '1' when (V_A_CTRL_INST_shadow /= R.A.CTRL.INST) else '0';
dfp_trap_vector(1967) <= '1' when (V_A_CTRL_PC_shadow /= RIN_D_PC_intermed_1) else '0';
dfp_trap_vector(1968) <= '1' when (V_A_CTRL_PC_shadow /= RIN_A_CTRL_PC_intermed_1) else '0';
dfp_trap_vector(1969) <= '1' when (V_A_CTRL_PC_shadow /= R.A.CTRL.PC) else '0';
dfp_trap_vector(1970) <= '1' when (V_A_CTRL_PC_shadow /= R.D.PC) else '0';
dfp_trap_vector(1971) <= '1' when (V_A_CTRL_PC_shadow /= V_D_PC_shadow_intermed_1) else '0';
dfp_trap_vector(1972) <= '1' when (V_A_CTRL_CNT_shadow /= RIN_D_CNT_intermed_1) else '0';
dfp_trap_vector(1973) <= '1' when (V_A_CTRL_CNT_shadow /= R.A.CTRL.CNT) else '0';
dfp_trap_vector(1974) <= '1' when (V_A_CTRL_CNT_shadow /= V_D_CNT_shadow_intermed_1) else '0';
dfp_trap_vector(1975) <= '1' when (V_A_CTRL_CNT_shadow /= R.D.CNT) else '0';
dfp_trap_vector(1976) <= '1' when (V_A_CTRL_CNT_shadow /= RIN_A_CTRL_CNT_intermed_1) else '0';
dfp_trap_vector(1977) <= '1' when (V_A_CTRL_CNT_shadow /= "00") else '0';
dfp_trap_vector(1978) <= '1' when (V_A_STEP_shadow /= R_D_ANNUL_intermed_1) else '0';
dfp_trap_vector(1979) <= '1' when (V_A_STEP_shadow /= RIN_D_STEP_intermed_1) else '0';
dfp_trap_vector(1980) <= '1' when (V_A_STEP_shadow /= V_D_ANNUL_shadow_intermed_2) else '0';
dfp_trap_vector(1981) <= '1' when (V_A_STEP_shadow /= R.A.STEP) else '0';
dfp_trap_vector(1982) <= '1' when (V_A_STEP_shadow /= DBGI_STEP_intermed_1) else '0';
dfp_trap_vector(1983) <= '1' when (V_A_STEP_shadow /= V_D_STEP_shadow_intermed_1) else '0';
dfp_trap_vector(1984) <= '1' when (V_A_STEP_shadow /= RIN_D_ANNUL_intermed_2) else '0';
dfp_trap_vector(1985) <= '1' when (V_A_STEP_shadow /= R.D.STEP) else '0';
dfp_trap_vector(1986) <= '1' when (V_A_STEP_shadow /= RIN_A_STEP_intermed_1) else '0';
dfp_trap_vector(1987) <= '1' when (V_D_STEP_shadow /= R.D.ANNUL) else '0';
dfp_trap_vector(1988) <= '1' when (V_D_STEP_shadow /= RIN_D_STEP_intermed_1) else '0';
dfp_trap_vector(1989) <= '1' when (V_D_STEP_shadow /= V_D_ANNUL_shadow_intermed_1) else '0';
dfp_trap_vector(1990) <= '1' when (V_D_STEP_shadow /= DBGI.STEP) else '0';
dfp_trap_vector(1991) <= '1' when (V_D_STEP_shadow /= RIN_D_ANNUL_intermed_1) else '0';
dfp_trap_vector(1992) <= '1' when (V_D_STEP_shadow /= R.D.STEP) else '0';
dfp_trap_vector(1993) <= '1' when (V_D_CNT_shadow /= RIN_D_CNT_intermed_1) else '0';
dfp_trap_vector(1994) <= '1' when (V_D_CNT_shadow /= R.D.CNT) else '0';
dfp_trap_vector(1995) <= '1' when (V_D_CNT_shadow /= "00") else '0';
dfp_trap_vector(1996) <= '1' when (V_F_PC_shadow /= EX_ADD_RES32DOWNTO3_shadow_intermed_1) else '0';
dfp_trap_vector(1997) <= '1' when (V_F_PC_shadow /= XC_TRAP_ADDRESS_shadow) else '0';
dfp_trap_vector(1998) <= '1' when (V_F_PC_shadow /= RIN_F_PC_intermed_1) else '0';
dfp_trap_vector(1999) <= '1' when (V_F_PC_shadow /= R.F.PC) else '0';
dfp_trap_vector(2000) <= '1' when (V_F_PC_shadow /= EX_JUMP_ADDRESS_shadow_intermed_1) else '0';
dfp_trap_vector(2001) <= '1' when (V_F_PC_shadow /= "000000000000000000000000000000") else '0';
dfp_trap_vector(2002) <= '1' when (V_F_BRANCH_shadow /= RIN_F_BRANCH_intermed_1) else '0';
dfp_trap_vector(2003) <= '1' when (V_F_BRANCH_shadow /= '1') else '0';
dfp_trap_vector(2004) <= '1' when (V_F_BRANCH_shadow /= '0') else '0';
dfp_trap_vector(2005) <= '1' when (V_F_BRANCH_shadow /= R.F.BRANCH) else '0';
dfp_trap_vector(2006) <= '1' when (V_F_PC31DOWNTO12_shadow /= R.F.PC ( 31 DOWNTO 12 )) else '0';
dfp_trap_vector(2007) <= '1' when (V_F_PC31DOWNTO12_shadow /= R_M_CTRL_PC31DOWNTO12_intermed_3) else '0';
dfp_trap_vector(2008) <= '1' when (V_F_PC31DOWNTO12_shadow /= V_D_PC31DOWNTO12_shadow_intermed_7) else '0';
dfp_trap_vector(2009) <= '1' when (V_F_PC31DOWNTO12_shadow /= V_A_CTRL_PC31DOWNTO12_shadow_intermed_6) else '0';
dfp_trap_vector(2010) <= '1' when (V_F_PC31DOWNTO12_shadow /= V_E_CTRL_PC31DOWNTO12_shadow_intermed_5) else '0';
dfp_trap_vector(2011) <= '1' when (V_F_PC31DOWNTO12_shadow /= EX_ADD_RES32DOWNTO330DOWNTO11_shadow_intermed_2) else '0';
dfp_trap_vector(2012) <= '1' when (V_F_PC31DOWNTO12_shadow /= RIN_F_PC31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(2013) <= '1' when (V_F_PC31DOWNTO12_shadow /= R_A_CTRL_PC31DOWNTO12_intermed_5) else '0';
dfp_trap_vector(2014) <= '1' when (V_F_PC31DOWNTO12_shadow /= R_E_CTRL_PC31DOWNTO12_intermed_4) else '0';
dfp_trap_vector(2015) <= '1' when (V_F_PC31DOWNTO12_shadow /= EX_JUMP_ADDRESS31DOWNTO12_shadow_intermed_2) else '0';
dfp_trap_vector(2016) <= '1' when (V_F_PC31DOWNTO12_shadow /= RIN_F_PC31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(2017) <= '1' when (V_F_PC31DOWNTO12_shadow /= RIN_A_CTRL_PC31DOWNTO12_intermed_6) else '0';
dfp_trap_vector(2018) <= '1' when (V_F_PC31DOWNTO12_shadow /= RIN_E_CTRL_PC31DOWNTO12_intermed_5) else '0';
dfp_trap_vector(2019) <= '1' when (V_F_PC31DOWNTO12_shadow /= V_F_PC31DOWNTO12_shadow_intermed_2) else '0';
dfp_trap_vector(2020) <= '1' when (V_F_PC31DOWNTO12_shadow /= IRIN_ADDR31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(2021) <= '1' when (V_F_PC31DOWNTO12_shadow /= V_X_CTRL_PC31DOWNTO12_shadow_intermed_3) else '0';
dfp_trap_vector(2022) <= '1' when (V_F_PC31DOWNTO12_shadow /= EX_ADD_RES32DOWNTO332DOWNTO13_shadow_intermed_2) else '0';
dfp_trap_vector(2023) <= '1' when (V_F_PC31DOWNTO12_shadow /= XC_TRAP_ADDRESS31DOWNTO12_shadow_intermed_1) else '0';
dfp_trap_vector(2024) <= '1' when (V_F_PC31DOWNTO12_shadow /= R_F_PC31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(2025) <= '1' when (V_F_PC31DOWNTO12_shadow /= RIN_M_CTRL_PC31DOWNTO12_intermed_4) else '0';
dfp_trap_vector(2026) <= '1' when (V_F_PC31DOWNTO12_shadow /= IR_ADDR31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(2027) <= '1' when (V_F_PC31DOWNTO12_shadow /= R_X_CTRL_PC31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(2028) <= '1' when (V_F_PC31DOWNTO12_shadow /= R_D_PC31DOWNTO12_intermed_6) else '0';
dfp_trap_vector(2029) <= '1' when (V_F_PC31DOWNTO12_shadow /= RIN_X_CTRL_PC31DOWNTO12_intermed_3) else '0';
dfp_trap_vector(2030) <= '1' when (V_F_PC31DOWNTO12_shadow /= RIN_D_PC31DOWNTO12_intermed_7) else '0';
dfp_trap_vector(2031) <= '1' when (V_F_PC31DOWNTO12_shadow /= VIR_ADDR31DOWNTO12_shadow_intermed_2) else '0';
dfp_trap_vector(2032) <= '1' when (V_F_PC31DOWNTO12_shadow /= V_M_CTRL_PC31DOWNTO12_shadow_intermed_4) else '0';
dfp_trap_vector(2033) <= '1' when (V_F_PC31DOWNTO2_shadow /= RIN_M_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2034) <= '1' when (V_F_PC31DOWNTO2_shadow /= V_D_PC31DOWNTO2_shadow_intermed_7) else '0';
dfp_trap_vector(2035) <= '1' when (V_F_PC31DOWNTO2_shadow /= RIN_D_PC31DOWNTO2_intermed_7) else '0';
dfp_trap_vector(2036) <= '1' when (V_F_PC31DOWNTO2_shadow /= EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_2) else '0';
dfp_trap_vector(2037) <= '1' when (V_F_PC31DOWNTO2_shadow /= V_F_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2038) <= '1' when (V_F_PC31DOWNTO2_shadow /= RIN_F_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2039) <= '1' when (V_F_PC31DOWNTO2_shadow /= RIN_X_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2040) <= '1' when (V_F_PC31DOWNTO2_shadow /= IRIN_ADDR31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2041) <= '1' when (V_F_PC31DOWNTO2_shadow /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_6) else '0';
dfp_trap_vector(2042) <= '1' when (V_F_PC31DOWNTO2_shadow(29 downto 2) /= X"0000001") else '0';
dfp_trap_vector(2043) <= '1' when (V_F_PC31DOWNTO2_shadow /= R_D_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(2044) <= '1' when (V_F_PC31DOWNTO2_shadow /= R.F.PC ( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(2045) <= '1' when (V_F_PC31DOWNTO2_shadow /= R_F_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2046) <= '1' when (V_F_PC31DOWNTO2_shadow /= VIR_ADDR31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2047) <= '1' when (V_F_PC31DOWNTO2_shadow /= R_M_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2048) <= '1' when (V_F_PC31DOWNTO2_shadow /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(2049) <= '1' when (V_F_PC31DOWNTO2_shadow /= RIN_A_CTRL_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(2050) <= '1' when (V_F_PC31DOWNTO2_shadow /= R_A_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2051) <= '1' when (V_F_PC31DOWNTO2_shadow /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(2052) <= '1' when (V_F_PC31DOWNTO2_shadow /= R_X_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2053) <= '1' when (V_F_PC31DOWNTO2_shadow /= XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(2054) <= '1' when (V_F_PC31DOWNTO2_shadow /= R_E_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2055) <= '1' when (V_F_PC31DOWNTO2_shadow /= EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2056) <= '1' when (V_F_PC31DOWNTO2_shadow /= RIN_F_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2057) <= '1' when (V_F_PC31DOWNTO2_shadow /= IR_ADDR31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2058) <= '1' when (V_F_PC31DOWNTO2_shadow /= RIN_E_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2059) <= '1' when (V_F_PC31DOWNTO2_shadow /= V_X_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(2060) <= '1' when (NPC31DOWNTO2_shadow /= RIN_M_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2061) <= '1' when (NPC31DOWNTO2_shadow /= V_D_PC31DOWNTO2_shadow_intermed_7) else '0';
dfp_trap_vector(2062) <= '1' when (NPC31DOWNTO2_shadow /= RIN_D_PC31DOWNTO2_intermed_7) else '0';
dfp_trap_vector(2063) <= '1' when (NPC31DOWNTO2_shadow /= EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_1) else '0';
dfp_trap_vector(2064) <= '1' when (NPC31DOWNTO2_shadow /= V_F_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(2065) <= '1' when (NPC31DOWNTO2_shadow /= RIN_F_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2066) <= '1' when (NPC31DOWNTO2_shadow /= RIN_X_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2067) <= '1' when (NPC31DOWNTO2_shadow /= IRIN_ADDR31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2068) <= '1' when (NPC31DOWNTO2_shadow /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_6) else '0';
dfp_trap_vector(2069) <= '1' when (NPC31DOWNTO2_shadow /= R_D_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(2070) <= '1' when (NPC31DOWNTO2_shadow /= R.F.PC( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(2071) <= '1' when (NPC31DOWNTO2_shadow /= VIR_ADDR31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2072) <= '1' when (NPC31DOWNTO2_shadow /= R_M_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2073) <= '1' when (NPC31DOWNTO2_shadow /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(2074) <= '1' when (NPC31DOWNTO2_shadow /= RIN_A_CTRL_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(2075) <= '1' when (NPC31DOWNTO2_shadow /= R_A_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2076) <= '1' when (NPC31DOWNTO2_shadow /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(2077) <= '1' when (NPC31DOWNTO2_shadow /= R_X_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2078) <= '1' when (NPC31DOWNTO2_shadow /= XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(2079) <= '1' when (NPC31DOWNTO2_shadow /= R_E_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2080) <= '1' when (NPC31DOWNTO2_shadow /= EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(2081) <= '1' when (NPC31DOWNTO2_shadow /= IR_ADDR31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2082) <= '1' when (NPC31DOWNTO2_shadow /= RIN_E_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2083) <= '1' when (NPC31DOWNTO2_shadow /= V_X_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(2084) <= '1' when (V_D_INST0_shadow /= RIN_D_INST0_intermed_1) else '0';
dfp_trap_vector(2085) <= '1' when (V_D_INST0_shadow /= R_D_INST0_intermed_1) else '0';
dfp_trap_vector(2086) <= '1' when (V_D_INST0_shadow /= R.D.INST ( 0 )) else '0';
dfp_trap_vector(2087) <= '1' when (V_D_INST0_shadow /= ICO.DATA ( 0 )) else '0';
dfp_trap_vector(2088) <= '1' when (V_D_INST0_shadow /= V_D_INST0_shadow_intermed_2) else '0';
dfp_trap_vector(2089) <= '1' when (V_D_INST0_shadow /= RIN_D_INST0_intermed_2) else '0';
dfp_trap_vector(2090) <= '1' when (V_D_INST1_shadow /= RIN_D_INST1_intermed_1) else '0';
dfp_trap_vector(2091) <= '1' when (V_D_INST1_shadow /= R_D_INST1_intermed_1) else '0';
dfp_trap_vector(2092) <= '1' when (V_D_INST1_shadow /= R.D.INST ( 1 )) else '0';
dfp_trap_vector(2093) <= '1' when (V_D_INST1_shadow /= ICO.DATA ( 1 )) else '0';
dfp_trap_vector(2094) <= '1' when (V_D_INST1_shadow /= V_D_INST1_shadow_intermed_2) else '0';
dfp_trap_vector(2095) <= '1' when (V_D_INST1_shadow /= RIN_D_INST1_intermed_2) else '0';
dfp_trap_vector(2096) <= '1' when (V_D_SET_shadow /= ICO.SET ( 0 DOWNTO 0 )) else '0';
dfp_trap_vector(2097) <= '1' when (V_D_SET_shadow /= R.D.SET) else '0';
dfp_trap_vector(2098) <= '1' when (V_D_SET_shadow /= RIN_D_SET_intermed_1) else '0';
dfp_trap_vector(2099) <= '1' when (V_D_MEXC_shadow /= ICO.MEXC) else '0';
dfp_trap_vector(2100) <= '1' when (V_D_MEXC_shadow /= R.D.MEXC) else '0';
dfp_trap_vector(2101) <= '1' when (V_D_MEXC_shadow /= RIN_D_MEXC_intermed_1) else '0';
dfp_trap_vector(2102) <= '1' when (EX_OP131_shadow /= RIN_X_DATA031_intermed_1) else '0';
dfp_trap_vector(2103) <= '1' when (EX_OP131_shadow /= RIN_E_OP131_intermed_1) else '0';
dfp_trap_vector(2104) <= '1' when (EX_OP131_shadow /= V_X_DATA031_shadow_intermed_1) else '0';
dfp_trap_vector(2105) <= '1' when (EX_OP131_shadow /= R.E.OP1( 31 )) else '0';
dfp_trap_vector(2106) <= '1' when (EX_OP131_shadow /= V_X_DATA031_shadow_intermed_2) else '0';
dfp_trap_vector(2107) <= '1' when (EX_OP131_shadow /= RIN_X_DATA031_intermed_2) else '0';
dfp_trap_vector(2108) <= '1' when (EX_OP131_shadow /= DCO_DATA031_intermed_1) else '0';
dfp_trap_vector(2109) <= '1' when (EX_OP131_shadow /= V_E_OP131_shadow_intermed_1) else '0';
dfp_trap_vector(2110) <= '1' when (EX_OP131_shadow /= R_X_DATA031_intermed_1) else '0';
dfp_trap_vector(2111) <= '1' when (EX_OP131_shadow /= R.X.DATA ( 0 )( 31 )) else '0';
dfp_trap_vector(2112) <= '1' when (EX_OP231_shadow /= RIN_X_DATA031_intermed_1) else '0';
dfp_trap_vector(2113) <= '1' when (EX_OP231_shadow /= V_X_DATA031_shadow_intermed_1) else '0';
dfp_trap_vector(2114) <= '1' when (EX_OP231_shadow /= V_X_DATA031_shadow_intermed_2) else '0';
dfp_trap_vector(2115) <= '1' when (EX_OP231_shadow /= RIN_X_DATA031_intermed_2) else '0';
dfp_trap_vector(2116) <= '1' when (EX_OP231_shadow /= DCO_DATA031_intermed_1) else '0';
dfp_trap_vector(2117) <= '1' when (EX_OP231_shadow /= RIN_E_OP231_intermed_1) else '0';
dfp_trap_vector(2118) <= '1' when (EX_OP231_shadow /= R_X_DATA031_intermed_1) else '0';
dfp_trap_vector(2119) <= '1' when (EX_OP231_shadow /= R.E.OP2( 31 )) else '0';
dfp_trap_vector(2120) <= '1' when (EX_OP231_shadow /= V_E_OP231_shadow_intermed_1) else '0';
dfp_trap_vector(2121) <= '1' when (EX_OP231_shadow /= R.X.DATA ( 0 )( 31 )) else '0';
dfp_trap_vector(2122) <= '1' when (VFPI_D_ANNUL_shadow /= R.D.ANNUL) else '0';
dfp_trap_vector(2123) <= '1' when (VFPI_D_ANNUL_shadow /= R.X.ANNUL_ALL) else '0';
dfp_trap_vector(2124) <= '1' when (VFPI_D_ANNUL_shadow /= '1') else '0';
dfp_trap_vector(2125) <= '1' when (VFPI_D_ANNUL_shadow /= '0') else '0';
dfp_trap_vector(2126) <= '1' when (VFPI_D_ANNUL_shadow /= V_D_ANNUL_shadow_intermed_1) else '0';
dfp_trap_vector(2127) <= '1' when (VFPI_D_ANNUL_shadow /= V_X_ANNUL_ALL_shadow) else '0';
dfp_trap_vector(2128) <= '1' when (VFPI_D_ANNUL_shadow /= RIN_X_ANNUL_ALL_intermed_1) else '0';
dfp_trap_vector(2129) <= '1' when (VFPI_D_ANNUL_shadow /= RIN_D_ANNUL_intermed_1) else '0';
dfp_trap_vector(2130) <= '1' when (VFPI_DBG_ENABLE_shadow /= '0') else '0';
dfp_trap_vector(2131) <= '1' when (VFPI_DBG_ENABLE_shadow /= DBGI.DENABLE) else '0';
dfp_trap_vector(2132) <= '1' when (EX_OP13_shadow /= V_X_DATA03_shadow_intermed_2) else '0';
dfp_trap_vector(2133) <= '1' when (EX_OP13_shadow /= V_X_DATA03_shadow_intermed_1) else '0';
dfp_trap_vector(2134) <= '1' when (EX_OP13_shadow /= DCO_DATA03_intermed_1) else '0';
dfp_trap_vector(2135) <= '1' when (EX_OP13_shadow /= RIN_X_DATA03_intermed_1) else '0';
dfp_trap_vector(2136) <= '1' when (EX_OP13_shadow /= R_X_DATA03_intermed_1) else '0';
dfp_trap_vector(2137) <= '1' when (EX_OP13_shadow /= RIN_X_DATA03_intermed_2) else '0';
dfp_trap_vector(2138) <= '1' when (EX_OP13_shadow /= RIN_E_OP13_intermed_1) else '0';
dfp_trap_vector(2139) <= '1' when (EX_OP13_shadow /= R.X.DATA ( 0 )( 3 )) else '0';
dfp_trap_vector(2140) <= '1' when (EX_OP13_shadow /= R.E.OP1( 3 )) else '0';
dfp_trap_vector(2141) <= '1' when (EX_OP13_shadow /= V_E_OP13_shadow_intermed_1) else '0';
dfp_trap_vector(2142) <= '1' when (EX_OP23_shadow /= V_X_DATA03_shadow_intermed_2) else '0';
dfp_trap_vector(2143) <= '1' when (EX_OP23_shadow /= V_X_DATA03_shadow_intermed_1) else '0';
dfp_trap_vector(2144) <= '1' when (EX_OP23_shadow /= DCO_DATA03_intermed_1) else '0';
dfp_trap_vector(2145) <= '1' when (EX_OP23_shadow /= R.E.OP2( 3 )) else '0';
dfp_trap_vector(2146) <= '1' when (EX_OP23_shadow /= RIN_X_DATA03_intermed_1) else '0';
dfp_trap_vector(2147) <= '1' when (EX_OP23_shadow /= R_X_DATA03_intermed_1) else '0';
dfp_trap_vector(2148) <= '1' when (EX_OP23_shadow /= RIN_X_DATA03_intermed_2) else '0';
dfp_trap_vector(2149) <= '1' when (EX_OP23_shadow /= RIN_E_OP23_intermed_1) else '0';
dfp_trap_vector(2150) <= '1' when (EX_OP23_shadow /= R.X.DATA ( 0 )( 3 )) else '0';
dfp_trap_vector(2151) <= '1' when (EX_OP23_shadow /= V_E_OP23_shadow_intermed_1) else '0';
dfp_trap_vector(2152) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= R_M_CTRL_PC31DOWNTO12_intermed_3) else '0';
dfp_trap_vector(2153) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= V_D_PC31DOWNTO12_shadow_intermed_7) else '0';
dfp_trap_vector(2154) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= V_A_CTRL_PC31DOWNTO12_shadow_intermed_6) else '0';
dfp_trap_vector(2155) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= V_E_CTRL_PC31DOWNTO12_shadow_intermed_5) else '0';
dfp_trap_vector(2156) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= EX_ADD_RES32DOWNTO330DOWNTO11_shadow_intermed_1) else '0';
dfp_trap_vector(2157) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= RIN_F_PC31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(2158) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= R_A_CTRL_PC31DOWNTO12_intermed_5) else '0';
dfp_trap_vector(2159) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= R_E_CTRL_PC31DOWNTO12_intermed_4) else '0';
dfp_trap_vector(2160) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= EX_JUMP_ADDRESS31DOWNTO12_shadow_intermed_1) else '0';
dfp_trap_vector(2161) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= RIN_A_CTRL_PC31DOWNTO12_intermed_6) else '0';
dfp_trap_vector(2162) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= RIN_E_CTRL_PC31DOWNTO12_intermed_5) else '0';
dfp_trap_vector(2163) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= V_F_PC31DOWNTO12_shadow_intermed_1) else '0';
dfp_trap_vector(2164) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= IRIN_ADDR31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(2165) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= V_X_CTRL_PC31DOWNTO12_shadow_intermed_3) else '0';
dfp_trap_vector(2166) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= EX_ADD_RES32DOWNTO332DOWNTO13_shadow_intermed_1) else '0';
dfp_trap_vector(2167) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= R.F.PC( 31 DOWNTO 12 )) else '0';
dfp_trap_vector(2168) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= RIN_M_CTRL_PC31DOWNTO12_intermed_4) else '0';
dfp_trap_vector(2169) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= IR_ADDR31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(2170) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= R_X_CTRL_PC31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(2171) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= R_D_PC31DOWNTO12_intermed_6) else '0';
dfp_trap_vector(2172) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= RIN_X_CTRL_PC31DOWNTO12_intermed_3) else '0';
dfp_trap_vector(2173) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= RIN_D_PC31DOWNTO12_intermed_7) else '0';
dfp_trap_vector(2174) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= VIR_ADDR31DOWNTO12_shadow_intermed_2) else '0';
dfp_trap_vector(2175) <= '1' when (XC_TRAP_ADDRESS31DOWNTO12_shadow /= V_M_CTRL_PC31DOWNTO12_shadow_intermed_4) else '0';
dfp_trap_vector(2176) <= '1' when (EX_JUMP_ADDRESS31DOWNTO12_shadow /= EX_ADD_RES32DOWNTO330DOWNTO11_shadow) else '0';
dfp_trap_vector(2177) <= '1' when (EX_JUMP_ADDRESS31DOWNTO12_shadow /= EX_ADD_RES32DOWNTO332DOWNTO13_shadow) else '0';
dfp_trap_vector(2178) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= RIN_M_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2179) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= V_D_PC31DOWNTO2_shadow_intermed_7) else '0';
dfp_trap_vector(2180) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= RIN_D_PC31DOWNTO2_intermed_7) else '0';
dfp_trap_vector(2181) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_1) else '0';
dfp_trap_vector(2182) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= V_F_PC31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(2183) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= RIN_F_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2184) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= RIN_X_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2185) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= IRIN_ADDR31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2186) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_6) else '0';
dfp_trap_vector(2187) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= R_D_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(2188) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= R.F.PC( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(2189) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= VIR_ADDR31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2190) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= R_M_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2191) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(2192) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= RIN_A_CTRL_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(2193) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= R_A_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2194) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(2195) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= R_X_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2196) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= R_E_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2197) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(2198) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= IR_ADDR31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2199) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= RIN_E_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2200) <= '1' when (XC_TRAP_ADDRESS31DOWNTO2_shadow /= V_X_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(2201) <= '1' when (V_F_PC31DOWNTO2_shadow /= RIN_M_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2202) <= '1' when (V_F_PC31DOWNTO2_shadow /= V_D_PC31DOWNTO2_shadow_intermed_7) else '0';
dfp_trap_vector(2203) <= '1' when (V_F_PC31DOWNTO2_shadow /= RIN_D_PC31DOWNTO2_intermed_7) else '0';
dfp_trap_vector(2204) <= '1' when (V_F_PC31DOWNTO2_shadow /= EX_ADD_RES32DOWNTO332DOWNTO3_shadow_intermed_1) else '0';
dfp_trap_vector(2205) <= '1' when (V_F_PC31DOWNTO2_shadow /= RIN_F_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2206) <= '1' when (V_F_PC31DOWNTO2_shadow /= RIN_X_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2207) <= '1' when (V_F_PC31DOWNTO2_shadow /= IRIN_ADDR31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2208) <= '1' when (V_F_PC31DOWNTO2_shadow /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_6) else '0';
dfp_trap_vector(2209) <= '1' when (V_F_PC31DOWNTO2_shadow /= R_D_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(2210) <= '1' when (V_F_PC31DOWNTO2_shadow /= R.F.PC( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(2211) <= '1' when (V_F_PC31DOWNTO2_shadow /= VIR_ADDR31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2212) <= '1' when (V_F_PC31DOWNTO2_shadow /= R_M_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2213) <= '1' when (V_F_PC31DOWNTO2_shadow /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(2214) <= '1' when (V_F_PC31DOWNTO2_shadow /= RIN_A_CTRL_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(2215) <= '1' when (V_F_PC31DOWNTO2_shadow /= R_A_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2216) <= '1' when (V_F_PC31DOWNTO2_shadow /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(2217) <= '1' when (V_F_PC31DOWNTO2_shadow /= R_X_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2218) <= '1' when (V_F_PC31DOWNTO2_shadow /= XC_TRAP_ADDRESS31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(2219) <= '1' when (V_F_PC31DOWNTO2_shadow /= R_E_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2220) <= '1' when (V_F_PC31DOWNTO2_shadow /= EX_JUMP_ADDRESS31DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(2221) <= '1' when (V_F_PC31DOWNTO2_shadow /= IR_ADDR31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2222) <= '1' when (V_F_PC31DOWNTO2_shadow /= RIN_E_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2223) <= '1' when (V_F_PC31DOWNTO2_shadow /= V_X_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(2224) <= '1' when (EX_OP231_shadow /= RIN_X_DATA031_intermed_1) else '0';
dfp_trap_vector(2225) <= '1' when (EX_OP231_shadow /= V_X_DATA031_shadow_intermed_1) else '0';
dfp_trap_vector(2226) <= '1' when (EX_OP231_shadow /= V_X_DATA031_shadow_intermed_2) else '0';
dfp_trap_vector(2227) <= '1' when (EX_OP231_shadow /= RIN_X_DATA031_intermed_2) else '0';
dfp_trap_vector(2228) <= '1' when (EX_OP231_shadow /= DCO_DATA031_intermed_1) else '0';
dfp_trap_vector(2229) <= '1' when (EX_OP231_shadow /= RIN_E_OP231_intermed_1) else '0';
dfp_trap_vector(2230) <= '1' when (EX_OP231_shadow /= R_X_DATA031_intermed_1) else '0';
dfp_trap_vector(2231) <= '1' when (EX_OP231_shadow /= R.E.OP2( 31 )) else '0';
dfp_trap_vector(2232) <= '1' when (EX_OP231_shadow /= V_E_OP231_shadow_intermed_1) else '0';
dfp_trap_vector(2233) <= '1' when (EX_OP231_shadow /= R.X.DATA ( 0 )( 31 )) else '0';
dfp_trap_vector(2234) <= '1' when (V_X_CTRL_RD7DOWNTO0_shadow /= V_M_CTRL_RD7DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(2235) <= '1' when (V_X_CTRL_RD7DOWNTO0_shadow /= V_E_CTRL_RD7DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(2236) <= '1' when (V_X_CTRL_RD7DOWNTO0_shadow /= R_E_CTRL_RD7DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2237) <= '1' when (V_X_CTRL_RD7DOWNTO0_shadow /= R.X.CTRL.RD ( 7 DOWNTO 0 )) else '0';
dfp_trap_vector(2238) <= '1' when (V_X_CTRL_RD7DOWNTO0_shadow /= V_A_CTRL_RD7DOWNTO0_shadow_intermed_4) else '0';
dfp_trap_vector(2239) <= '1' when (V_X_CTRL_RD7DOWNTO0_shadow /= RIN_A_CTRL_RD7DOWNTO0_intermed_4) else '0';
dfp_trap_vector(2240) <= '1' when (V_X_CTRL_RD7DOWNTO0_shadow /= R_M_CTRL_RD7DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2241) <= '1' when (V_X_CTRL_RD7DOWNTO0_shadow /= R_A_CTRL_RD7DOWNTO0_intermed_3) else '0';
dfp_trap_vector(2242) <= '1' when (V_X_CTRL_RD7DOWNTO0_shadow /= RIN_E_CTRL_RD7DOWNTO0_intermed_3) else '0';
dfp_trap_vector(2243) <= '1' when (V_X_CTRL_RD7DOWNTO0_shadow /= RIN_X_CTRL_RD7DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2244) <= '1' when (V_X_CTRL_RD7DOWNTO0_shadow /= RIN_M_CTRL_RD7DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2245) <= '1' when (V_X_CTRL_TRAP_shadow /= RIN_X_CTRL_TRAP_intermed_1) else '0';
dfp_trap_vector(2246) <= '1' when (V_X_CTRL_TRAP_shadow /= V_A_CTRL_TRAP_shadow_intermed_4) else '0';
dfp_trap_vector(2247) <= '1' when (V_X_CTRL_TRAP_shadow /= ICO_MEXC_intermed_5) else '0';
dfp_trap_vector(2248) <= '1' when (V_X_CTRL_TRAP_shadow /= R_E_CTRL_TRAP_intermed_2) else '0';
dfp_trap_vector(2249) <= '1' when (V_X_CTRL_TRAP_shadow /= RIN_A_CTRL_TRAP_intermed_4) else '0';
dfp_trap_vector(2250) <= '1' when (V_X_CTRL_TRAP_shadow /= V_E_CTRL_TRAP_shadow_intermed_3) else '0';
dfp_trap_vector(2251) <= '1' when (V_X_CTRL_TRAP_shadow /= RIN_E_CTRL_TRAP_intermed_3) else '0';
dfp_trap_vector(2252) <= '1' when (V_X_CTRL_TRAP_shadow /= R_D_MEXC_intermed_4) else '0';
dfp_trap_vector(2253) <= '1' when (V_X_CTRL_TRAP_shadow /= R.X.CTRL.TRAP) else '0';
dfp_trap_vector(2254) <= '1' when (V_X_CTRL_TRAP_shadow /= V_M_CTRL_TRAP_shadow_intermed_2) else '0';
dfp_trap_vector(2255) <= '1' when (V_X_CTRL_TRAP_shadow /= V_D_MEXC_shadow_intermed_5) else '0';
dfp_trap_vector(2256) <= '1' when (V_X_CTRL_TRAP_shadow /= R_A_CTRL_TRAP_intermed_3) else '0';
dfp_trap_vector(2257) <= '1' when (V_X_CTRL_TRAP_shadow /= RIN_M_CTRL_TRAP_intermed_2) else '0';
dfp_trap_vector(2258) <= '1' when (V_X_CTRL_TRAP_shadow /= R_M_CTRL_TRAP_intermed_1) else '0';
dfp_trap_vector(2259) <= '1' when (V_X_CTRL_TRAP_shadow /= RIN_D_MEXC_intermed_5) else '0';
dfp_trap_vector(2260) <= '1' when (V_X_RESULT6DOWNTO0_shadow /= RIN_X_RESULT6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2261) <= '1' when (V_X_RESULT6DOWNTO0_shadow /= R.X.RESULT ( 6 DOWNTO 0 )) else '0';
dfp_trap_vector(2262) <= '1' when (V_X_RESULT6DOWNTO0_shadow /= V_X_RESULT6DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(2263) <= '1' when (V_X_RESULT6DOWNTO0_shadow /= RIN_X_RESULT6DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2264) <= '1' when (V_X_RESULT6DOWNTO0_shadow /= R_X_RESULT6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2265) <= '1' when (V_X_CTRL_PC_shadow /= RIN_D_PC_intermed_5) else '0';
dfp_trap_vector(2266) <= '1' when (V_X_CTRL_PC_shadow /= RIN_A_CTRL_PC_intermed_4) else '0';
dfp_trap_vector(2267) <= '1' when (V_X_CTRL_PC_shadow /= R_A_CTRL_PC_intermed_3) else '0';
dfp_trap_vector(2268) <= '1' when (V_X_CTRL_PC_shadow /= V_E_CTRL_PC_shadow_intermed_3) else '0';
dfp_trap_vector(2269) <= '1' when (V_X_CTRL_PC_shadow /= R_M_CTRL_PC_intermed_1) else '0';
dfp_trap_vector(2270) <= '1' when (V_X_CTRL_PC_shadow /= R.X.CTRL.PC) else '0';
dfp_trap_vector(2271) <= '1' when (V_X_CTRL_PC_shadow /= R_E_CTRL_PC_intermed_2) else '0';
dfp_trap_vector(2272) <= '1' when (V_X_CTRL_PC_shadow /= RIN_M_CTRL_PC_intermed_2) else '0';
dfp_trap_vector(2273) <= '1' when (V_X_CTRL_PC_shadow /= V_M_CTRL_PC_shadow_intermed_2) else '0';
dfp_trap_vector(2274) <= '1' when (V_X_CTRL_PC_shadow /= V_A_CTRL_PC_shadow_intermed_4) else '0';
dfp_trap_vector(2275) <= '1' when (V_X_CTRL_PC_shadow /= R_D_PC_intermed_4) else '0';
dfp_trap_vector(2276) <= '1' when (V_X_CTRL_PC_shadow /= RIN_E_CTRL_PC_intermed_3) else '0';
dfp_trap_vector(2277) <= '1' when (V_X_CTRL_PC_shadow /= RIN_X_CTRL_PC_intermed_1) else '0';
dfp_trap_vector(2278) <= '1' when (V_X_CTRL_PC_shadow /= V_D_PC_shadow_intermed_5) else '0';
dfp_trap_vector(2279) <= '1' when (V_X_CTRL_WREG_shadow /= RIN_A_CTRL_ANNUL_intermed_5) else '0';
dfp_trap_vector(2280) <= '1' when (V_X_CTRL_WREG_shadow /= R.X.CTRL.WREG) else '0';
dfp_trap_vector(2281) <= '1' when (V_X_CTRL_WREG_shadow /= R_A_CTRL_ANNUL_intermed_4) else '0';
dfp_trap_vector(2282) <= '1' when (V_X_CTRL_WREG_shadow /= R_X_ANNUL_ALL_intermed_4) else '0';
dfp_trap_vector(2283) <= '1' when (V_X_CTRL_WREG_shadow /= RIN_X_CTRL_WREG_intermed_1) else '0';
dfp_trap_vector(2284) <= '1' when (V_X_CTRL_WREG_shadow /= '1') else '0';
dfp_trap_vector(2285) <= '1' when (V_X_CTRL_WREG_shadow /= '0') else '0';
dfp_trap_vector(2286) <= '1' when (V_X_CTRL_WREG_shadow /= RIN_M_CTRL_WREG_intermed_2) else '0';
dfp_trap_vector(2287) <= '1' when (V_X_CTRL_WREG_shadow /= RIN_A_CTRL_WREG_intermed_4) else '0';
dfp_trap_vector(2288) <= '1' when (V_X_CTRL_WREG_shadow /= V_A_CTRL_WREG_shadow_intermed_4) else '0';
dfp_trap_vector(2289) <= '1' when (V_X_CTRL_WREG_shadow /= R_A_CTRL_WREG_intermed_3) else '0';
dfp_trap_vector(2290) <= '1' when (V_X_CTRL_WREG_shadow /= V_X_ANNUL_ALL_shadow_intermed_4) else '0';
dfp_trap_vector(2291) <= '1' when (V_X_CTRL_WREG_shadow /= R_M_CTRL_WREG_intermed_1) else '0';
dfp_trap_vector(2292) <= '1' when (V_X_CTRL_WREG_shadow /= RIN_X_ANNUL_ALL_intermed_5) else '0';
dfp_trap_vector(2293) <= '1' when (V_X_CTRL_WREG_shadow /= V_M_CTRL_WREG_shadow_intermed_2) else '0';
dfp_trap_vector(2294) <= '1' when (V_X_CTRL_WREG_shadow /= R_E_CTRL_WREG_intermed_2) else '0';
dfp_trap_vector(2295) <= '1' when (V_X_CTRL_WREG_shadow /= V_A_CTRL_ANNUL_shadow_intermed_4) else '0';
dfp_trap_vector(2296) <= '1' when (V_X_CTRL_WREG_shadow /= RIN_E_CTRL_WREG_intermed_3) else '0';
dfp_trap_vector(2297) <= '1' when (V_X_CTRL_WREG_shadow /= V_E_CTRL_WREG_shadow_intermed_3) else '0';
dfp_trap_vector(2298) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= RIN_M_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2299) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2300) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= R_E_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2301) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= V_D_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(2302) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= RIN_D_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2303) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= RIN_E_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2304) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= RIN_A_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2305) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= RIN_X_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2306) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= RIN_X_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2307) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= RIN_M_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2308) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= R.X.CTRL.PC ( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(2309) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(2310) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= R_D_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2311) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= R_M_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2312) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= R_M_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2313) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(2314) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= RIN_A_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2315) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= R_A_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2316) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(2317) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= R_A_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2318) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= R_X_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2319) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(2320) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= R_E_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2321) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= RIN_E_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2322) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= V_X_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2323) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(2324) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= RIN_M_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2325) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= V_D_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(2326) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= RIN_D_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2327) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= RIN_X_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2328) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(2329) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= R_D_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2330) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= R_M_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2331) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(2332) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= RIN_A_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2333) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= R_A_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2334) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2335) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= R.X.CTRL.PC( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(2336) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= R_E_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2337) <= '1' when (V_X_CTRL_PC31DOWNTO2_shadow /= RIN_E_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2338) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= V_X_CTRL_TT3DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(2339) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= R_M_CTRL_TT3DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2340) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(2341) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= R_X_RESULT6DOWNTO03DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2342) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= R_A_CTRL_TT3DOWNTO0_intermed_4) else '0';
dfp_trap_vector(2343) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= RIN_A_CTRL_TT3DOWNTO0_intermed_5) else '0';
dfp_trap_vector(2344) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= V_A_CTRL_TT3DOWNTO0_shadow_intermed_5) else '0';
dfp_trap_vector(2345) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= RIN_W_S_TT3DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2346) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= R_E_CTRL_TT3DOWNTO0_intermed_3) else '0';
dfp_trap_vector(2347) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= RIN_W_S_TT3DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2348) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= RIN_M_CTRL_TT3DOWNTO0_intermed_3) else '0';
dfp_trap_vector(2349) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= V_M_CTRL_TT3DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(2350) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_3) else '0';
dfp_trap_vector(2351) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2352) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= R_W_S_TT3DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2353) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= R_X_RESULT6DOWNTO03DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2354) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(2355) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= V_E_CTRL_TT3DOWNTO0_shadow_intermed_4) else '0';
dfp_trap_vector(2356) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= RIN_X_CTRL_TT3DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2357) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= V_W_S_TT3DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(2358) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= R_X_CTRL_TT3DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2359) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= RIN_E_CTRL_TT3DOWNTO0_intermed_4) else '0';
dfp_trap_vector(2360) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= R.W.S.TT ( 3 DOWNTO 0 )) else '0';
dfp_trap_vector(2361) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= XC_VECTT3DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(2362) <= '1' when (V_M_RESULT1DOWNTO0_shadow /= V_M_RESULT1DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(2363) <= '1' when (V_M_RESULT1DOWNTO0_shadow /= R.M.RESULT ( 1 DOWNTO 0 )) else '0';
dfp_trap_vector(2364) <= '1' when (V_M_RESULT1DOWNTO0_shadow /= RIN_M_RESULT1DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2365) <= '1' when (V_M_RESULT1DOWNTO0_shadow /= R_M_RESULT1DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2366) <= '1' when (V_M_RESULT1DOWNTO0_shadow /= RIN_M_RESULT1DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2367) <= '1' when (V_X_DATA031_shadow /= RIN_X_DATA031_intermed_2) else '0';
dfp_trap_vector(2368) <= '1' when (V_X_DATA031_shadow /= V_X_DATA031_shadow_intermed_2) else '0';
dfp_trap_vector(2369) <= '1' when (V_X_DATA031_shadow /= V_X_DATA031_shadow_intermed_3) else '0';
dfp_trap_vector(2370) <= '1' when (V_X_DATA031_shadow /= RIN_X_DATA031_intermed_3) else '0';
dfp_trap_vector(2371) <= '1' when (V_X_DATA031_shadow /= DCO_DATA031_intermed_1) else '0';
dfp_trap_vector(2372) <= '1' when (V_X_DATA031_shadow /= R.X.DATA ( 0 ) ( 31 )) else '0';
dfp_trap_vector(2373) <= '1' when (V_X_DATA031_shadow /= RIN_X_DATA031_intermed_1) else '0';
dfp_trap_vector(2374) <= '1' when (V_X_DATA031_shadow /= R_X_DATA031_intermed_2) else '0';
dfp_trap_vector(2375) <= '1' when (V_X_DATA031_shadow /= R_X_DATA031_intermed_1) else '0';
dfp_trap_vector(2376) <= '1' when (V_X_DATA031_shadow /= RIN_X_DATA031_intermed_1) else '0';
dfp_trap_vector(2377) <= '1' when (V_X_DATA031_shadow /= V_X_DATA031_shadow_intermed_2) else '0';
dfp_trap_vector(2378) <= '1' when (V_X_DATA031_shadow /= RIN_X_DATA031_intermed_2) else '0';
dfp_trap_vector(2379) <= '1' when (V_X_DATA031_shadow /= DCO_DATA031_intermed_1) else '0';
dfp_trap_vector(2380) <= '1' when (V_X_DATA031_shadow /= R_X_DATA031_intermed_1) else '0';
dfp_trap_vector(2381) <= '1' when (V_X_DATA031_shadow /= R.X.DATA ( 0 )( 31 )) else '0';
dfp_trap_vector(2382) <= '1' when (V_E_CTRL_INST19_shadow /= V_A_CTRL_INST19_shadow_intermed_3) else '0';
dfp_trap_vector(2383) <= '1' when (V_E_CTRL_INST19_shadow /= V_E_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(2384) <= '1' when (V_E_CTRL_INST19_shadow /= RIN_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(2385) <= '1' when (V_E_CTRL_INST19_shadow /= RIN_A_CTRL_INST19_intermed_3) else '0';
dfp_trap_vector(2386) <= '1' when (V_E_CTRL_INST19_shadow /= RIN_E_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(2387) <= '1' when (V_E_CTRL_INST19_shadow /= R.E.CTRL.INST ( 19 )) else '0';
dfp_trap_vector(2388) <= '1' when (V_E_CTRL_INST19_shadow /= RIN_E_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(2389) <= '1' when (V_E_CTRL_INST19_shadow /= DE_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(2390) <= '1' when (V_E_CTRL_INST19_shadow /= R_E_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(2391) <= '1' when (V_E_CTRL_INST19_shadow /= R_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(2392) <= '1' when (V_E_CTRL_INST19_shadow /= R_A_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(2393) <= '1' when (V_E_CTRL_INST19_shadow /= V_A_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(2394) <= '1' when (V_E_CTRL_INST20_shadow /= R.E.CTRL.INST ( 20 )) else '0';
dfp_trap_vector(2395) <= '1' when (V_E_CTRL_INST20_shadow /= RIN_A_CTRL_INST20_intermed_2) else '0';
dfp_trap_vector(2396) <= '1' when (V_E_CTRL_INST20_shadow /= R_A_CTRL_INST20_intermed_1) else '0';
dfp_trap_vector(2397) <= '1' when (V_E_CTRL_INST20_shadow /= RIN_A_CTRL_INST20_intermed_3) else '0';
dfp_trap_vector(2398) <= '1' when (V_E_CTRL_INST20_shadow /= V_E_CTRL_INST20_shadow_intermed_2) else '0';
dfp_trap_vector(2399) <= '1' when (V_E_CTRL_INST20_shadow /= V_A_CTRL_INST20_shadow_intermed_3) else '0';
dfp_trap_vector(2400) <= '1' when (V_E_CTRL_INST20_shadow /= RIN_E_CTRL_INST20_intermed_2) else '0';
dfp_trap_vector(2401) <= '1' when (V_E_CTRL_INST20_shadow /= V_A_CTRL_INST20_shadow_intermed_2) else '0';
dfp_trap_vector(2402) <= '1' when (V_E_CTRL_INST20_shadow /= RIN_E_CTRL_INST20_intermed_1) else '0';
dfp_trap_vector(2403) <= '1' when (V_E_CTRL_INST20_shadow /= R_E_CTRL_INST20_intermed_1) else '0';
dfp_trap_vector(2404) <= '1' when (V_E_CTRL_INST20_shadow /= DE_INST20_shadow_intermed_2) else '0';
dfp_trap_vector(2405) <= '1' when (V_E_CTRL_INST20_shadow /= R_A_CTRL_INST20_intermed_2) else '0';
dfp_trap_vector(2406) <= '1' when (V_X_DATA00_shadow /= V_X_DATA00_shadow_intermed_2) else '0';
dfp_trap_vector(2407) <= '1' when (V_X_DATA00_shadow /= R.X.DATA ( 0 ) ( 0 )) else '0';
dfp_trap_vector(2408) <= '1' when (V_X_DATA00_shadow /= RIN_X_DATA00_intermed_1) else '0';
dfp_trap_vector(2409) <= '1' when (V_X_DATA00_shadow /= R_X_DATA00_intermed_2) else '0';
dfp_trap_vector(2410) <= '1' when (V_X_DATA00_shadow /= RIN_X_DATA00_intermed_2) else '0';
dfp_trap_vector(2411) <= '1' when (V_X_DATA00_shadow /= DCO_DATA00_intermed_1) else '0';
dfp_trap_vector(2412) <= '1' when (V_X_DATA00_shadow /= V_X_DATA00_shadow_intermed_3) else '0';
dfp_trap_vector(2413) <= '1' when (V_X_DATA00_shadow /= R_X_DATA00_intermed_1) else '0';
dfp_trap_vector(2414) <= '1' when (V_X_DATA00_shadow /= RIN_X_DATA00_intermed_3) else '0';
dfp_trap_vector(2415) <= '1' when (V_X_DATA00_shadow /= R_X_DATA00_intermed_1) else '0';
dfp_trap_vector(2416) <= '1' when (V_X_DATA00_shadow /= RIN_X_DATA00_intermed_1) else '0';
dfp_trap_vector(2417) <= '1' when (V_X_DATA00_shadow /= DCO_DATA00_intermed_1) else '0';
dfp_trap_vector(2418) <= '1' when (V_X_DATA00_shadow /= V_X_DATA00_shadow_intermed_2) else '0';
dfp_trap_vector(2419) <= '1' when (V_X_DATA00_shadow /= R.X.DATA ( 0 )( 0 )) else '0';
dfp_trap_vector(2420) <= '1' when (V_X_DATA00_shadow /= RIN_X_DATA00_intermed_2) else '0';
dfp_trap_vector(2421) <= '1' when (V_X_DATA04DOWNTO0_shadow /= RIN_X_DATA04DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2422) <= '1' when (V_X_DATA04DOWNTO0_shadow /= R_X_DATA04DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2423) <= '1' when (V_X_DATA04DOWNTO0_shadow /= R_X_DATA04DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2424) <= '1' when (V_X_DATA04DOWNTO0_shadow /= RIN_X_DATA04DOWNTO0_intermed_3) else '0';
dfp_trap_vector(2425) <= '1' when (V_X_DATA04DOWNTO0_shadow /= R.X.DATA ( 0 ) ( 4 DOWNTO 0 )) else '0';
dfp_trap_vector(2426) <= '1' when (V_X_DATA04DOWNTO0_shadow /= V_X_DATA04DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(2427) <= '1' when (V_X_DATA04DOWNTO0_shadow /= V_X_DATA04DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(2428) <= '1' when (V_X_DATA04DOWNTO0_shadow /= RIN_X_DATA04DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2429) <= '1' when (V_X_DATA04DOWNTO0_shadow /= DCO_DATA04DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2430) <= '1' when (V_X_DATA04DOWNTO0_shadow /= R_X_DATA04DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2431) <= '1' when (V_X_DATA04DOWNTO0_shadow /= R.X.DATA ( 0 )( 4 DOWNTO 0 )) else '0';
dfp_trap_vector(2432) <= '1' when (V_X_DATA04DOWNTO0_shadow /= RIN_X_DATA04DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2433) <= '1' when (V_X_DATA04DOWNTO0_shadow /= V_X_DATA04DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(2434) <= '1' when (V_X_DATA04DOWNTO0_shadow /= DCO_DATA04DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2435) <= '1' when (V_X_DATA04DOWNTO0_shadow /= RIN_X_DATA04DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2436) <= '1' when (V_D_PC31DOWNTO2_shadow /= V_D_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2437) <= '1' when (V_D_PC31DOWNTO2_shadow /= RIN_D_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2438) <= '1' when (V_D_PC31DOWNTO2_shadow /= R_D_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2439) <= '1' when (V_D_PC31DOWNTO2_shadow /= R.D.PC ( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(2440) <= '1' when (V_D_PC31DOWNTO2_shadow /= RIN_D_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2441) <= '1' when (V_E_CTRL_INST24_shadow /= R_A_CTRL_INST24_intermed_2) else '0';
dfp_trap_vector(2442) <= '1' when (V_E_CTRL_INST24_shadow /= RIN_E_CTRL_INST24_intermed_2) else '0';
dfp_trap_vector(2443) <= '1' when (V_E_CTRL_INST24_shadow /= RIN_A_CTRL_INST24_intermed_3) else '0';
dfp_trap_vector(2444) <= '1' when (V_E_CTRL_INST24_shadow /= R_E_CTRL_INST24_intermed_1) else '0';
dfp_trap_vector(2445) <= '1' when (V_E_CTRL_INST24_shadow /= R_A_CTRL_INST24_intermed_1) else '0';
dfp_trap_vector(2446) <= '1' when (V_E_CTRL_INST24_shadow /= R.E.CTRL.INST ( 24 )) else '0';
dfp_trap_vector(2447) <= '1' when (V_E_CTRL_INST24_shadow /= V_A_CTRL_INST24_shadow_intermed_3) else '0';
dfp_trap_vector(2448) <= '1' when (V_E_CTRL_INST24_shadow /= V_E_CTRL_INST24_shadow_intermed_2) else '0';
dfp_trap_vector(2449) <= '1' when (V_E_CTRL_INST24_shadow /= DE_INST24_shadow_intermed_2) else '0';
dfp_trap_vector(2450) <= '1' when (V_E_CTRL_INST24_shadow /= RIN_A_CTRL_INST24_intermed_2) else '0';
dfp_trap_vector(2451) <= '1' when (V_E_CTRL_INST24_shadow /= V_A_CTRL_INST24_shadow_intermed_2) else '0';
dfp_trap_vector(2452) <= '1' when (V_E_CTRL_INST24_shadow /= RIN_E_CTRL_INST24_intermed_1) else '0';
dfp_trap_vector(2453) <= '1' when (V_A_CTRL_INST19_shadow /= V_A_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(2454) <= '1' when (V_A_CTRL_INST19_shadow /= RIN_A_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(2455) <= '1' when (V_A_CTRL_INST19_shadow /= RIN_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(2456) <= '1' when (V_A_CTRL_INST19_shadow /= DE_INST19_shadow_intermed_1) else '0';
dfp_trap_vector(2457) <= '1' when (V_A_CTRL_INST19_shadow /= R_A_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(2458) <= '1' when (V_A_CTRL_INST19_shadow /= R.A.CTRL.INST ( 19 )) else '0';
dfp_trap_vector(2459) <= '1' when (V_M_Y31_shadow /= RIN_M_Y31_intermed_1) else '0';
dfp_trap_vector(2460) <= '1' when (V_M_Y31_shadow /= V_M_Y31_shadow_intermed_2) else '0';
dfp_trap_vector(2461) <= '1' when (V_M_Y31_shadow /= RIN_M_Y31_intermed_2) else '0';
dfp_trap_vector(2462) <= '1' when (V_M_Y31_shadow /= R_M_Y31_intermed_1) else '0';
dfp_trap_vector(2463) <= '1' when (V_M_Y31_shadow /= R.M.Y ( 31 )) else '0';
dfp_trap_vector(2464) <= '1' when (VDSU_CRDY2_shadow /= DSUIN_CRDY2_intermed_1) else '0';
dfp_trap_vector(2465) <= '1' when (VDSU_CRDY2_shadow /= DSUR.CRDY ( 2 )) else '0';
dfp_trap_vector(2466) <= '1' when (VDSU_CRDY2_shadow /= VDSU_CRDY2_shadow_intermed_2) else '0';
dfp_trap_vector(2467) <= '1' when (VDSU_CRDY2_shadow /= DSUIN_CRDY2_intermed_2) else '0';
dfp_trap_vector(2468) <= '1' when (VDSU_CRDY2_shadow /= DSUR_CRDY2_intermed_1) else '0';
dfp_trap_vector(2469) <= '1' when (V_A_CTRL_PC31DOWNTO2_shadow /= V_D_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2470) <= '1' when (V_A_CTRL_PC31DOWNTO2_shadow /= RIN_D_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2471) <= '1' when (V_A_CTRL_PC31DOWNTO2_shadow /= RIN_A_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2472) <= '1' when (V_A_CTRL_PC31DOWNTO2_shadow /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2473) <= '1' when (V_A_CTRL_PC31DOWNTO2_shadow /= R_D_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2474) <= '1' when (V_A_CTRL_PC31DOWNTO2_shadow /= RIN_A_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2475) <= '1' when (V_A_CTRL_PC31DOWNTO2_shadow /= R_A_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2476) <= '1' when (V_A_CTRL_PC31DOWNTO2_shadow /= R.A.CTRL.PC ( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(2477) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= R.E.CTRL.PC ( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(2478) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= V_D_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(2479) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= RIN_D_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2480) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= RIN_E_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2481) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= RIN_A_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2482) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(2483) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= R_D_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2484) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2485) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= RIN_A_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2486) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= R_A_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2487) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= R_A_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2488) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2489) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= R_E_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2490) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= RIN_E_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2491) <= '1' when (V_E_CTRL_INST_shadow /= R.E.CTRL.INST) else '0';
dfp_trap_vector(2492) <= '1' when (V_E_CTRL_INST_shadow /= DE_INST_shadow_intermed_2) else '0';
dfp_trap_vector(2493) <= '1' when (V_E_CTRL_INST_shadow /= V_A_CTRL_INST_shadow_intermed_2) else '0';
dfp_trap_vector(2494) <= '1' when (V_E_CTRL_INST_shadow /= RIN_A_CTRL_INST_intermed_2) else '0';
dfp_trap_vector(2495) <= '1' when (V_E_CTRL_INST_shadow /= RIN_E_CTRL_INST_intermed_1) else '0';
dfp_trap_vector(2496) <= '1' when (V_E_CTRL_INST_shadow /= R_A_CTRL_INST_intermed_1) else '0';
dfp_trap_vector(2497) <= '1' when (V_E_CTRL_CNT_shadow /= RIN_D_CNT_intermed_3) else '0';
dfp_trap_vector(2498) <= '1' when (V_E_CTRL_CNT_shadow /= V_A_CTRL_CNT_shadow_intermed_2) else '0';
dfp_trap_vector(2499) <= '1' when (V_E_CTRL_CNT_shadow /= R_A_CTRL_CNT_intermed_1) else '0';
dfp_trap_vector(2500) <= '1' when (V_E_CTRL_CNT_shadow /= V_D_CNT_shadow_intermed_3) else '0';
dfp_trap_vector(2501) <= '1' when (V_E_CTRL_CNT_shadow /= R_D_CNT_intermed_2) else '0';
dfp_trap_vector(2502) <= '1' when (V_E_CTRL_CNT_shadow /= R.E.CTRL.CNT) else '0';
dfp_trap_vector(2503) <= '1' when (V_E_CTRL_CNT_shadow /= RIN_A_CTRL_CNT_intermed_2) else '0';
dfp_trap_vector(2504) <= '1' when (V_E_CTRL_CNT_shadow /= "00") else '0';
dfp_trap_vector(2505) <= '1' when (V_E_CTRL_CNT_shadow /= RIN_E_CTRL_CNT_intermed_1) else '0';
dfp_trap_vector(2506) <= '1' when (V_E_CTRL_TRAP_shadow /= V_A_CTRL_TRAP_shadow_intermed_2) else '0';
dfp_trap_vector(2507) <= '1' when (V_E_CTRL_TRAP_shadow /= ICO_MEXC_intermed_3) else '0';
dfp_trap_vector(2508) <= '1' when (V_E_CTRL_TRAP_shadow /= R.E.CTRL.TRAP) else '0';
dfp_trap_vector(2509) <= '1' when (V_E_CTRL_TRAP_shadow /= RIN_A_CTRL_TRAP_intermed_2) else '0';
dfp_trap_vector(2510) <= '1' when (V_E_CTRL_TRAP_shadow /= RIN_E_CTRL_TRAP_intermed_1) else '0';
dfp_trap_vector(2511) <= '1' when (V_E_CTRL_TRAP_shadow /= R_D_MEXC_intermed_2) else '0';
dfp_trap_vector(2512) <= '1' when (V_E_CTRL_TRAP_shadow /= V_D_MEXC_shadow_intermed_3) else '0';
dfp_trap_vector(2513) <= '1' when (V_E_CTRL_TRAP_shadow /= R_A_CTRL_TRAP_intermed_1) else '0';
dfp_trap_vector(2514) <= '1' when (V_E_CTRL_TRAP_shadow /= RIN_D_MEXC_intermed_3) else '0';
dfp_trap_vector(2515) <= '1' when (V_E_CTRL_PV_shadow /= R.E.CTRL.PV) else '0';
dfp_trap_vector(2516) <= '1' when (V_E_CTRL_PV_shadow /= R_A_CTRL_PV_intermed_1) else '0';
dfp_trap_vector(2517) <= '1' when (V_E_CTRL_PV_shadow /= RIN_E_CTRL_PV_intermed_1) else '0';
dfp_trap_vector(2518) <= '1' when (V_E_CTRL_PV_shadow /= V_A_CTRL_PV_shadow_intermed_2) else '0';
dfp_trap_vector(2519) <= '1' when (V_E_CTRL_PV_shadow /= RIN_A_CTRL_PV_intermed_2) else '0';
dfp_trap_vector(2520) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= RIN_M_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2521) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= R_E_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2522) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= V_D_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(2523) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= RIN_D_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2524) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= RIN_E_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2525) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= RIN_A_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2526) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= RIN_M_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2527) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(2528) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= R_D_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2529) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= R.M.CTRL.PC ( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(2530) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= R_M_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2531) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(2532) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= RIN_A_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2533) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= R_A_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2534) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2535) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= R_A_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2536) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(2537) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= R_E_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2538) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= RIN_E_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2539) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2540) <= '1' when (V_M_CTRL_INST_shadow /= R_E_CTRL_INST_intermed_1) else '0';
dfp_trap_vector(2541) <= '1' when (V_M_CTRL_INST_shadow /= R.M.CTRL.INST) else '0';
dfp_trap_vector(2542) <= '1' when (V_M_CTRL_INST_shadow /= DE_INST_shadow_intermed_3) else '0';
dfp_trap_vector(2543) <= '1' when (V_M_CTRL_INST_shadow /= V_A_CTRL_INST_shadow_intermed_3) else '0';
dfp_trap_vector(2544) <= '1' when (V_M_CTRL_INST_shadow /= V_E_CTRL_INST_shadow_intermed_2) else '0';
dfp_trap_vector(2545) <= '1' when (V_M_CTRL_INST_shadow /= RIN_A_CTRL_INST_intermed_3) else '0';
dfp_trap_vector(2546) <= '1' when (V_M_CTRL_INST_shadow /= RIN_M_CTRL_INST_intermed_1) else '0';
dfp_trap_vector(2547) <= '1' when (V_M_CTRL_INST_shadow /= RIN_E_CTRL_INST_intermed_2) else '0';
dfp_trap_vector(2548) <= '1' when (V_M_CTRL_INST_shadow /= R_A_CTRL_INST_intermed_2) else '0';
dfp_trap_vector(2549) <= '1' when (V_M_CTRL_CNT_shadow /= V_E_CTRL_CNT_shadow_intermed_2) else '0';
dfp_trap_vector(2550) <= '1' when (V_M_CTRL_CNT_shadow /= RIN_D_CNT_intermed_4) else '0';
dfp_trap_vector(2551) <= '1' when (V_M_CTRL_CNT_shadow /= R.M.CTRL.CNT) else '0';
dfp_trap_vector(2552) <= '1' when (V_M_CTRL_CNT_shadow /= V_A_CTRL_CNT_shadow_intermed_3) else '0';
dfp_trap_vector(2553) <= '1' when (V_M_CTRL_CNT_shadow /= R_A_CTRL_CNT_intermed_2) else '0';
dfp_trap_vector(2554) <= '1' when (V_M_CTRL_CNT_shadow /= V_D_CNT_shadow_intermed_4) else '0';
dfp_trap_vector(2555) <= '1' when (V_M_CTRL_CNT_shadow /= R_D_CNT_intermed_3) else '0';
dfp_trap_vector(2556) <= '1' when (V_M_CTRL_CNT_shadow /= R_E_CTRL_CNT_intermed_1) else '0';
dfp_trap_vector(2557) <= '1' when (V_M_CTRL_CNT_shadow /= RIN_A_CTRL_CNT_intermed_3) else '0';
dfp_trap_vector(2558) <= '1' when (V_M_CTRL_CNT_shadow /= RIN_M_CTRL_CNT_intermed_1) else '0';
dfp_trap_vector(2559) <= '1' when (V_M_CTRL_CNT_shadow /= "00") else '0';
dfp_trap_vector(2560) <= '1' when (V_M_CTRL_CNT_shadow /= RIN_E_CTRL_CNT_intermed_2) else '0';
dfp_trap_vector(2561) <= '1' when (V_M_CTRL_TRAP_shadow /= V_A_CTRL_TRAP_shadow_intermed_3) else '0';
dfp_trap_vector(2562) <= '1' when (V_M_CTRL_TRAP_shadow /= ICO_MEXC_intermed_4) else '0';
dfp_trap_vector(2563) <= '1' when (V_M_CTRL_TRAP_shadow /= R_E_CTRL_TRAP_intermed_1) else '0';
dfp_trap_vector(2564) <= '1' when (V_M_CTRL_TRAP_shadow /= RIN_A_CTRL_TRAP_intermed_3) else '0';
dfp_trap_vector(2565) <= '1' when (V_M_CTRL_TRAP_shadow /= V_E_CTRL_TRAP_shadow_intermed_2) else '0';
dfp_trap_vector(2566) <= '1' when (V_M_CTRL_TRAP_shadow /= RIN_E_CTRL_TRAP_intermed_2) else '0';
dfp_trap_vector(2567) <= '1' when (V_M_CTRL_TRAP_shadow /= R_D_MEXC_intermed_3) else '0';
dfp_trap_vector(2568) <= '1' when (V_M_CTRL_TRAP_shadow /= V_D_MEXC_shadow_intermed_4) else '0';
dfp_trap_vector(2569) <= '1' when (V_M_CTRL_TRAP_shadow /= R_A_CTRL_TRAP_intermed_2) else '0';
dfp_trap_vector(2570) <= '1' when (V_M_CTRL_TRAP_shadow /= RIN_M_CTRL_TRAP_intermed_1) else '0';
dfp_trap_vector(2571) <= '1' when (V_M_CTRL_TRAP_shadow /= R.M.CTRL.TRAP) else '0';
dfp_trap_vector(2572) <= '1' when (V_M_CTRL_TRAP_shadow /= RIN_D_MEXC_intermed_4) else '0';
dfp_trap_vector(2573) <= '1' when (V_M_CTRL_PV_shadow /= V_E_CTRL_PV_shadow_intermed_2) else '0';
dfp_trap_vector(2574) <= '1' when (V_M_CTRL_PV_shadow /= R.M.CTRL.PV) else '0';
dfp_trap_vector(2575) <= '1' when (V_M_CTRL_PV_shadow /= R_E_CTRL_PV_intermed_1) else '0';
dfp_trap_vector(2576) <= '1' when (V_M_CTRL_PV_shadow /= R_A_CTRL_PV_intermed_2) else '0';
dfp_trap_vector(2577) <= '1' when (V_M_CTRL_PV_shadow /= RIN_E_CTRL_PV_intermed_2) else '0';
dfp_trap_vector(2578) <= '1' when (V_M_CTRL_PV_shadow /= RIN_M_CTRL_PV_intermed_1) else '0';
dfp_trap_vector(2579) <= '1' when (V_M_CTRL_PV_shadow /= V_A_CTRL_PV_shadow_intermed_3) else '0';
dfp_trap_vector(2580) <= '1' when (V_M_CTRL_PV_shadow /= RIN_A_CTRL_PV_intermed_3) else '0';
dfp_trap_vector(2581) <= '1' when (V_X_CTRL_INST_shadow /= R_E_CTRL_INST_intermed_2) else '0';
dfp_trap_vector(2582) <= '1' when (V_X_CTRL_INST_shadow /= R_M_CTRL_INST_intermed_1) else '0';
dfp_trap_vector(2583) <= '1' when (V_X_CTRL_INST_shadow /= DE_INST_shadow_intermed_4) else '0';
dfp_trap_vector(2584) <= '1' when (V_X_CTRL_INST_shadow /= V_A_CTRL_INST_shadow_intermed_4) else '0';
dfp_trap_vector(2585) <= '1' when (V_X_CTRL_INST_shadow /= V_E_CTRL_INST_shadow_intermed_3) else '0';
dfp_trap_vector(2586) <= '1' when (V_X_CTRL_INST_shadow /= R.X.CTRL.INST) else '0';
dfp_trap_vector(2587) <= '1' when (V_X_CTRL_INST_shadow /= RIN_X_CTRL_INST_intermed_1) else '0';
dfp_trap_vector(2588) <= '1' when (V_X_CTRL_INST_shadow /= RIN_A_CTRL_INST_intermed_4) else '0';
dfp_trap_vector(2589) <= '1' when (V_X_CTRL_INST_shadow /= RIN_M_CTRL_INST_intermed_2) else '0';
dfp_trap_vector(2590) <= '1' when (V_X_CTRL_INST_shadow /= RIN_E_CTRL_INST_intermed_3) else '0';
dfp_trap_vector(2591) <= '1' when (V_X_CTRL_INST_shadow /= V_M_CTRL_INST_shadow_intermed_2) else '0';
dfp_trap_vector(2592) <= '1' when (V_X_CTRL_INST_shadow /= R_A_CTRL_INST_intermed_3) else '0';
dfp_trap_vector(2593) <= '1' when (V_X_CTRL_CNT_shadow /= V_E_CTRL_CNT_shadow_intermed_3) else '0';
dfp_trap_vector(2594) <= '1' when (V_X_CTRL_CNT_shadow /= R.X.CTRL.CNT) else '0';
dfp_trap_vector(2595) <= '1' when (V_X_CTRL_CNT_shadow /= RIN_D_CNT_intermed_5) else '0';
dfp_trap_vector(2596) <= '1' when (V_X_CTRL_CNT_shadow /= R_M_CTRL_CNT_intermed_1) else '0';
dfp_trap_vector(2597) <= '1' when (V_X_CTRL_CNT_shadow /= V_A_CTRL_CNT_shadow_intermed_4) else '0';
dfp_trap_vector(2598) <= '1' when (V_X_CTRL_CNT_shadow /= R_A_CTRL_CNT_intermed_3) else '0';
dfp_trap_vector(2599) <= '1' when (V_X_CTRL_CNT_shadow /= V_D_CNT_shadow_intermed_5) else '0';
dfp_trap_vector(2600) <= '1' when (V_X_CTRL_CNT_shadow /= R_D_CNT_intermed_4) else '0';
dfp_trap_vector(2601) <= '1' when (V_X_CTRL_CNT_shadow /= R_E_CTRL_CNT_intermed_2) else '0';
dfp_trap_vector(2602) <= '1' when (V_X_CTRL_CNT_shadow /= RIN_X_CTRL_CNT_intermed_1) else '0';
dfp_trap_vector(2603) <= '1' when (V_X_CTRL_CNT_shadow /= RIN_A_CTRL_CNT_intermed_4) else '0';
dfp_trap_vector(2604) <= '1' when (V_X_CTRL_CNT_shadow /= RIN_M_CTRL_CNT_intermed_2) else '0';
dfp_trap_vector(2605) <= '1' when (V_X_CTRL_CNT_shadow /= "00") else '0';
dfp_trap_vector(2606) <= '1' when (V_X_CTRL_CNT_shadow /= RIN_E_CTRL_CNT_intermed_3) else '0';
dfp_trap_vector(2607) <= '1' when (V_X_CTRL_CNT_shadow /= V_M_CTRL_CNT_shadow_intermed_2) else '0';
dfp_trap_vector(2608) <= '1' when (V_X_CTRL_PV_shadow /= V_E_CTRL_PV_shadow_intermed_3) else '0';
dfp_trap_vector(2609) <= '1' when (V_X_CTRL_PV_shadow /= R_M_CTRL_PV_intermed_1) else '0';
dfp_trap_vector(2610) <= '1' when (V_X_CTRL_PV_shadow /= R_E_CTRL_PV_intermed_2) else '0';
dfp_trap_vector(2611) <= '1' when (V_X_CTRL_PV_shadow /= R_A_CTRL_PV_intermed_3) else '0';
dfp_trap_vector(2612) <= '1' when (V_X_CTRL_PV_shadow /= RIN_E_CTRL_PV_intermed_3) else '0';
dfp_trap_vector(2613) <= '1' when (V_X_CTRL_PV_shadow /= R.X.CTRL.PV) else '0';
dfp_trap_vector(2614) <= '1' when (V_X_CTRL_PV_shadow /= RIN_X_CTRL_PV_intermed_1) else '0';
dfp_trap_vector(2615) <= '1' when (V_X_CTRL_PV_shadow /= RIN_M_CTRL_PV_intermed_2) else '0';
dfp_trap_vector(2616) <= '1' when (V_X_CTRL_PV_shadow /= V_A_CTRL_PV_shadow_intermed_4) else '0';
dfp_trap_vector(2617) <= '1' when (V_X_CTRL_PV_shadow /= V_M_CTRL_PV_shadow_intermed_2) else '0';
dfp_trap_vector(2618) <= '1' when (V_X_CTRL_PV_shadow /= RIN_A_CTRL_PV_intermed_4) else '0';
dfp_trap_vector(2619) <= '1' when (V_E_CTRL_INST19_shadow /= V_A_CTRL_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(2620) <= '1' when (V_E_CTRL_INST19_shadow /= RIN_A_CTRL_INST19_intermed_2) else '0';
dfp_trap_vector(2621) <= '1' when (V_E_CTRL_INST19_shadow /= RIN_E_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(2622) <= '1' when (V_E_CTRL_INST19_shadow /= DE_INST19_shadow_intermed_2) else '0';
dfp_trap_vector(2623) <= '1' when (V_E_CTRL_INST19_shadow /= R.E.CTRL.INST( 19 )) else '0';
dfp_trap_vector(2624) <= '1' when (V_E_CTRL_INST19_shadow /= R_A_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(2625) <= '1' when (V_E_CTRL_INST20_shadow /= RIN_A_CTRL_INST20_intermed_2) else '0';
dfp_trap_vector(2626) <= '1' when (V_E_CTRL_INST20_shadow /= V_A_CTRL_INST20_shadow_intermed_2) else '0';
dfp_trap_vector(2627) <= '1' when (V_E_CTRL_INST20_shadow /= RIN_E_CTRL_INST20_intermed_1) else '0';
dfp_trap_vector(2628) <= '1' when (V_E_CTRL_INST20_shadow /= R.E.CTRL.INST( 20 )) else '0';
dfp_trap_vector(2629) <= '1' when (V_E_CTRL_INST20_shadow /= DE_INST20_shadow_intermed_2) else '0';
dfp_trap_vector(2630) <= '1' when (V_E_CTRL_INST20_shadow /= R_A_CTRL_INST20_intermed_1) else '0';
dfp_trap_vector(2631) <= '1' when (V_E_CTRL_INST24_shadow /= R_A_CTRL_INST24_intermed_1) else '0';
dfp_trap_vector(2632) <= '1' when (V_E_CTRL_INST24_shadow /= RIN_A_CTRL_INST24_intermed_2) else '0';
dfp_trap_vector(2633) <= '1' when (V_E_CTRL_INST24_shadow /= RIN_E_CTRL_INST24_intermed_1) else '0';
dfp_trap_vector(2634) <= '1' when (V_E_CTRL_INST24_shadow /= R.E.CTRL.INST( 24 )) else '0';
dfp_trap_vector(2635) <= '1' when (V_E_CTRL_INST24_shadow /= V_A_CTRL_INST24_shadow_intermed_2) else '0';
dfp_trap_vector(2636) <= '1' when (V_E_CTRL_INST24_shadow /= DE_INST24_shadow_intermed_2) else '0';
dfp_trap_vector(2637) <= '1' when (V_A_CTRL_INST19_shadow /= RIN_A_CTRL_INST19_intermed_1) else '0';
dfp_trap_vector(2638) <= '1' when (V_A_CTRL_INST19_shadow /= DE_INST19_shadow_intermed_1) else '0';
dfp_trap_vector(2639) <= '1' when (V_A_CTRL_INST19_shadow /= R.A.CTRL.INST( 19 )) else '0';
dfp_trap_vector(2640) <= '1' when (V_F_PC31DOWNTO4_shadow /= V_X_CTRL_PC31DOWNTO4_shadow_intermed_3) else '0';
dfp_trap_vector(2641) <= '1' when (V_F_PC31DOWNTO4_shadow /= IR_ADDR31DOWNTO4_intermed_1) else '0';
dfp_trap_vector(2642) <= '1' when (V_F_PC31DOWNTO4_shadow /= R.F.PC( 31 DOWNTO 4 )) else '0';
dfp_trap_vector(2643) <= '1' when (V_F_PC31DOWNTO4_shadow /= VIR_ADDR31DOWNTO4_shadow_intermed_2) else '0';
dfp_trap_vector(2644) <= '1' when (V_F_PC31DOWNTO4_shadow /= RIN_F_PC31DOWNTO4_intermed_1) else '0';
dfp_trap_vector(2645) <= '1' when (V_F_PC31DOWNTO4_shadow /= RIN_A_CTRL_PC31DOWNTO4_intermed_6) else '0';
dfp_trap_vector(2646) <= '1' when (V_F_PC31DOWNTO4_shadow /= R_A_CTRL_PC31DOWNTO4_intermed_5) else '0';
dfp_trap_vector(2647) <= '1' when (V_F_PC31DOWNTO4_shadow /= R_D_PC31DOWNTO4_intermed_6) else '0';
dfp_trap_vector(2648) <= '1' when (V_F_PC31DOWNTO4_shadow /= RIN_X_CTRL_PC31DOWNTO4_intermed_3) else '0';
dfp_trap_vector(2649) <= '1' when (V_F_PC31DOWNTO4_shadow /= EX_ADD_RES32DOWNTO332DOWNTO5_shadow_intermed_1) else '0';
dfp_trap_vector(2650) <= '1' when (V_F_PC31DOWNTO4_shadow /= V_D_PC31DOWNTO4_shadow_intermed_7) else '0';
dfp_trap_vector(2651) <= '1' when (V_F_PC31DOWNTO4_shadow /= V_E_CTRL_PC31DOWNTO4_shadow_intermed_5) else '0';
dfp_trap_vector(2652) <= '1' when (V_F_PC31DOWNTO4_shadow /= RIN_M_CTRL_PC31DOWNTO4_intermed_4) else '0';
dfp_trap_vector(2653) <= '1' when (V_F_PC31DOWNTO4_shadow /= R_X_CTRL_PC31DOWNTO4_intermed_2) else '0';
dfp_trap_vector(2654) <= '1' when (V_F_PC31DOWNTO4_shadow /= IRIN_ADDR31DOWNTO4_intermed_2) else '0';
dfp_trap_vector(2655) <= '1' when (V_F_PC31DOWNTO4_shadow /= V_M_CTRL_PC31DOWNTO4_shadow_intermed_4) else '0';
dfp_trap_vector(2656) <= '1' when (V_F_PC31DOWNTO4_shadow /= R_M_CTRL_PC31DOWNTO4_intermed_3) else '0';
dfp_trap_vector(2657) <= '1' when (V_F_PC31DOWNTO4_shadow /= XC_TRAP_ADDRESS31DOWNTO4_shadow_intermed_1) else '0';
dfp_trap_vector(2658) <= '1' when (V_F_PC31DOWNTO4_shadow /= RIN_D_PC31DOWNTO4_intermed_7) else '0';
dfp_trap_vector(2659) <= '1' when (V_F_PC31DOWNTO4_shadow /= RIN_E_CTRL_PC31DOWNTO4_intermed_5) else '0';
dfp_trap_vector(2660) <= '1' when (V_F_PC31DOWNTO4_shadow /= EX_JUMP_ADDRESS31DOWNTO4_shadow_intermed_1) else '0';
dfp_trap_vector(2661) <= '1' when (V_F_PC31DOWNTO4_shadow /= V_A_CTRL_PC31DOWNTO4_shadow_intermed_6) else '0';
dfp_trap_vector(2662) <= '1' when (V_F_PC31DOWNTO4_shadow /= R_E_CTRL_PC31DOWNTO4_intermed_4) else '0';
dfp_trap_vector(2663) <= '1' when (VIR_ADDR31DOWNTO4_shadow /= V_X_CTRL_PC31DOWNTO4_shadow_intermed_2) else '0';
dfp_trap_vector(2664) <= '1' when (VIR_ADDR31DOWNTO4_shadow /= IR.ADDR( 31 DOWNTO 4 )) else '0';
dfp_trap_vector(2665) <= '1' when (VIR_ADDR31DOWNTO4_shadow /= RIN_A_CTRL_PC31DOWNTO4_intermed_5) else '0';
dfp_trap_vector(2666) <= '1' when (VIR_ADDR31DOWNTO4_shadow /= R_A_CTRL_PC31DOWNTO4_intermed_4) else '0';
dfp_trap_vector(2667) <= '1' when (VIR_ADDR31DOWNTO4_shadow /= R_D_PC31DOWNTO4_intermed_5) else '0';
dfp_trap_vector(2668) <= '1' when (VIR_ADDR31DOWNTO4_shadow /= RIN_X_CTRL_PC31DOWNTO4_intermed_2) else '0';
dfp_trap_vector(2669) <= '1' when (VIR_ADDR31DOWNTO4_shadow /= V_D_PC31DOWNTO4_shadow_intermed_6) else '0';
dfp_trap_vector(2670) <= '1' when (VIR_ADDR31DOWNTO4_shadow /= V_E_CTRL_PC31DOWNTO4_shadow_intermed_4) else '0';
dfp_trap_vector(2671) <= '1' when (VIR_ADDR31DOWNTO4_shadow /= RIN_M_CTRL_PC31DOWNTO4_intermed_3) else '0';
dfp_trap_vector(2672) <= '1' when (VIR_ADDR31DOWNTO4_shadow /= R_X_CTRL_PC31DOWNTO4_intermed_1) else '0';
dfp_trap_vector(2673) <= '1' when (VIR_ADDR31DOWNTO4_shadow /= IRIN_ADDR31DOWNTO4_intermed_1) else '0';
dfp_trap_vector(2674) <= '1' when (VIR_ADDR31DOWNTO4_shadow /= V_M_CTRL_PC31DOWNTO4_shadow_intermed_3) else '0';
dfp_trap_vector(2675) <= '1' when (VIR_ADDR31DOWNTO4_shadow /= R_M_CTRL_PC31DOWNTO4_intermed_2) else '0';
dfp_trap_vector(2676) <= '1' when (VIR_ADDR31DOWNTO4_shadow /= RIN_D_PC31DOWNTO4_intermed_6) else '0';
dfp_trap_vector(2677) <= '1' when (VIR_ADDR31DOWNTO4_shadow /= RIN_E_CTRL_PC31DOWNTO4_intermed_4) else '0';
dfp_trap_vector(2678) <= '1' when (VIR_ADDR31DOWNTO4_shadow /= V_A_CTRL_PC31DOWNTO4_shadow_intermed_5) else '0';
dfp_trap_vector(2679) <= '1' when (VIR_ADDR31DOWNTO4_shadow /= R_E_CTRL_PC31DOWNTO4_intermed_3) else '0';
dfp_trap_vector(2680) <= '1' when (V_F_PC3DOWNTO2_shadow /= R_D_PC3DOWNTO2_intermed_6) else '0';
dfp_trap_vector(2681) <= '1' when (V_F_PC3DOWNTO2_shadow /= V_D_PC3DOWNTO2_shadow_intermed_7) else '0';
dfp_trap_vector(2682) <= '1' when (V_F_PC3DOWNTO2_shadow /= VIR_ADDR3DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2683) <= '1' when (V_F_PC3DOWNTO2_shadow /= RIN_D_PC3DOWNTO2_intermed_7) else '0';
dfp_trap_vector(2684) <= '1' when (V_F_PC3DOWNTO2_shadow /= R_M_CTRL_PC3DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2685) <= '1' when (V_F_PC3DOWNTO2_shadow /= R_E_CTRL_PC3DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2686) <= '1' when (V_F_PC3DOWNTO2_shadow /= V_E_CTRL_PC3DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(2687) <= '1' when (V_F_PC3DOWNTO2_shadow /= RIN_X_CTRL_PC3DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2688) <= '1' when (V_F_PC3DOWNTO2_shadow /= R_A_CTRL_PC3DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2689) <= '1' when (V_F_PC3DOWNTO2_shadow /= R.F.PC( 3 DOWNTO 2 )) else '0';
dfp_trap_vector(2690) <= '1' when (V_F_PC3DOWNTO2_shadow /= V_X_CTRL_PC3DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(2691) <= '1' when (V_F_PC3DOWNTO2_shadow /= RIN_M_CTRL_PC3DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2692) <= '1' when (V_F_PC3DOWNTO2_shadow /= IRIN_ADDR3DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2693) <= '1' when (V_F_PC3DOWNTO2_shadow /= EX_JUMP_ADDRESS3DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(2694) <= '1' when (V_F_PC3DOWNTO2_shadow /= EX_ADD_RES32DOWNTO34DOWNTO3_shadow_intermed_1) else '0';
dfp_trap_vector(2695) <= '1' when (V_F_PC3DOWNTO2_shadow /= RIN_A_CTRL_PC3DOWNTO2_intermed_6) else '0';
dfp_trap_vector(2696) <= '1' when (V_F_PC3DOWNTO2_shadow /= XC_TRAP_ADDRESS3DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(2697) <= '1' when (V_F_PC3DOWNTO2_shadow /= V_A_CTRL_PC3DOWNTO2_shadow_intermed_6) else '0';
dfp_trap_vector(2698) <= '1' when (V_F_PC3DOWNTO2_shadow /= IR_ADDR3DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2699) <= '1' when (V_F_PC3DOWNTO2_shadow /= V_M_CTRL_PC3DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(2700) <= '1' when (V_F_PC3DOWNTO2_shadow /= R_X_CTRL_PC3DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2701) <= '1' when (V_F_PC3DOWNTO2_shadow /= RIN_E_CTRL_PC3DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2702) <= '1' when (V_F_PC3DOWNTO2_shadow /= RIN_F_PC3DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2703) <= '1' when (VIR_ADDR3DOWNTO2_shadow /= R_D_PC3DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2704) <= '1' when (VIR_ADDR3DOWNTO2_shadow /= V_D_PC3DOWNTO2_shadow_intermed_6) else '0';
dfp_trap_vector(2705) <= '1' when (VIR_ADDR3DOWNTO2_shadow /= RIN_D_PC3DOWNTO2_intermed_6) else '0';
dfp_trap_vector(2706) <= '1' when (VIR_ADDR3DOWNTO2_shadow /= R_M_CTRL_PC3DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2707) <= '1' when (VIR_ADDR3DOWNTO2_shadow /= R_E_CTRL_PC3DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2708) <= '1' when (VIR_ADDR3DOWNTO2_shadow /= V_E_CTRL_PC3DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(2709) <= '1' when (VIR_ADDR3DOWNTO2_shadow /= RIN_X_CTRL_PC3DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2710) <= '1' when (VIR_ADDR3DOWNTO2_shadow /= R_A_CTRL_PC3DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2711) <= '1' when (VIR_ADDR3DOWNTO2_shadow /= V_X_CTRL_PC3DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2712) <= '1' when (VIR_ADDR3DOWNTO2_shadow /= RIN_M_CTRL_PC3DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2713) <= '1' when (VIR_ADDR3DOWNTO2_shadow /= IRIN_ADDR3DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2714) <= '1' when (VIR_ADDR3DOWNTO2_shadow /= RIN_A_CTRL_PC3DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2715) <= '1' when (VIR_ADDR3DOWNTO2_shadow /= V_A_CTRL_PC3DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(2716) <= '1' when (VIR_ADDR3DOWNTO2_shadow /= IR.ADDR( 3 DOWNTO 2 )) else '0';
dfp_trap_vector(2717) <= '1' when (VIR_ADDR3DOWNTO2_shadow /= V_M_CTRL_PC3DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(2718) <= '1' when (VIR_ADDR3DOWNTO2_shadow /= R_X_CTRL_PC3DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2719) <= '1' when (VIR_ADDR3DOWNTO2_shadow /= RIN_E_CTRL_PC3DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2720) <= '1' when (V_X_CTRL_RD6DOWNTO0_shadow /= RIN_E_CTRL_RD6DOWNTO0_intermed_3) else '0';
dfp_trap_vector(2721) <= '1' when (V_X_CTRL_RD6DOWNTO0_shadow /= RIN_M_CTRL_RD6DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2722) <= '1' when (V_X_CTRL_RD6DOWNTO0_shadow /= RIN_X_CTRL_RD6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2723) <= '1' when (V_X_CTRL_RD6DOWNTO0_shadow /= R.X.CTRL.RD( 6 DOWNTO 0 )) else '0';
dfp_trap_vector(2724) <= '1' when (V_X_CTRL_RD6DOWNTO0_shadow /= V_M_CTRL_RD6DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(2725) <= '1' when (V_X_CTRL_RD6DOWNTO0_shadow /= R_E_CTRL_RD6DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2726) <= '1' when (V_X_CTRL_RD6DOWNTO0_shadow /= V_E_CTRL_RD6DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(2727) <= '1' when (V_X_CTRL_RD6DOWNTO0_shadow /= V_A_CTRL_RD6DOWNTO0_shadow_intermed_4) else '0';
dfp_trap_vector(2728) <= '1' when (V_X_CTRL_RD6DOWNTO0_shadow /= R_A_CTRL_RD6DOWNTO0_intermed_3) else '0';
dfp_trap_vector(2729) <= '1' when (V_X_CTRL_RD6DOWNTO0_shadow /= RIN_A_CTRL_RD6DOWNTO0_intermed_4) else '0';
dfp_trap_vector(2730) <= '1' when (V_X_CTRL_RD6DOWNTO0_shadow /= R_M_CTRL_RD6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2731) <= '1' when (V_M_CTRL_TT_shadow /= V_E_CTRL_TT_shadow_intermed_2) else '0';
dfp_trap_vector(2732) <= '1' when (V_M_CTRL_TT_shadow /= RIN_A_CTRL_TT_intermed_3) else '0';
dfp_trap_vector(2733) <= '1' when (V_M_CTRL_TT_shadow /= R_A_CTRL_TT_intermed_2) else '0';
dfp_trap_vector(2734) <= '1' when (V_M_CTRL_TT_shadow /= R.M.CTRL.TT) else '0';
dfp_trap_vector(2735) <= '1' when (V_M_CTRL_TT_shadow /= "000000") else '0';
dfp_trap_vector(2736) <= '1' when (V_M_CTRL_TT_shadow /= R_E_CTRL_TT_intermed_1) else '0';
dfp_trap_vector(2737) <= '1' when (V_M_CTRL_TT_shadow /= RIN_M_CTRL_TT_intermed_1) else '0';
dfp_trap_vector(2738) <= '1' when (V_M_CTRL_TT_shadow /= RIN_E_CTRL_TT_intermed_2) else '0';
dfp_trap_vector(2739) <= '1' when (V_M_CTRL_TT_shadow /= V_A_CTRL_TT_shadow_intermed_3) else '0';
dfp_trap_vector(2740) <= '1' when (V_E_CTRL_LD_shadow /= R_A_CTRL_LD_intermed_1) else '0';
dfp_trap_vector(2741) <= '1' when (V_E_CTRL_LD_shadow /= RIN_A_CTRL_LD_intermed_2) else '0';
dfp_trap_vector(2742) <= '1' when (V_E_CTRL_LD_shadow /= R.E.CTRL.LD) else '0';
dfp_trap_vector(2743) <= '1' when (V_E_CTRL_LD_shadow /= RIN_E_CTRL_LD_intermed_1) else '0';
dfp_trap_vector(2744) <= '1' when (V_E_CTRL_LD_shadow /= V_A_CTRL_LD_shadow_intermed_2) else '0';
dfp_trap_vector(2745) <= '1' when (V_F_PC31DOWNTO12_shadow /= R_M_CTRL_PC31DOWNTO12_intermed_3) else '0';
dfp_trap_vector(2746) <= '1' when (V_F_PC31DOWNTO12_shadow /= V_D_PC31DOWNTO12_shadow_intermed_7) else '0';
dfp_trap_vector(2747) <= '1' when (V_F_PC31DOWNTO12_shadow /= V_A_CTRL_PC31DOWNTO12_shadow_intermed_6) else '0';
dfp_trap_vector(2748) <= '1' when (V_F_PC31DOWNTO12_shadow /= V_E_CTRL_PC31DOWNTO12_shadow_intermed_5) else '0';
dfp_trap_vector(2749) <= '1' when (V_F_PC31DOWNTO12_shadow /= EX_ADD_RES32DOWNTO330DOWNTO11_shadow_intermed_1) else '0';
dfp_trap_vector(2750) <= '1' when (V_F_PC31DOWNTO12_shadow /= RIN_F_PC31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(2751) <= '1' when (V_F_PC31DOWNTO12_shadow /= R_A_CTRL_PC31DOWNTO12_intermed_5) else '0';
dfp_trap_vector(2752) <= '1' when (V_F_PC31DOWNTO12_shadow /= R_E_CTRL_PC31DOWNTO12_intermed_4) else '0';
dfp_trap_vector(2753) <= '1' when (V_F_PC31DOWNTO12_shadow /= EX_JUMP_ADDRESS31DOWNTO12_shadow_intermed_1) else '0';
dfp_trap_vector(2754) <= '1' when (V_F_PC31DOWNTO12_shadow /= RIN_A_CTRL_PC31DOWNTO12_intermed_6) else '0';
dfp_trap_vector(2755) <= '1' when (V_F_PC31DOWNTO12_shadow /= RIN_E_CTRL_PC31DOWNTO12_intermed_5) else '0';
dfp_trap_vector(2756) <= '1' when (V_F_PC31DOWNTO12_shadow /= IRIN_ADDR31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(2757) <= '1' when (V_F_PC31DOWNTO12_shadow /= V_X_CTRL_PC31DOWNTO12_shadow_intermed_3) else '0';
dfp_trap_vector(2758) <= '1' when (V_F_PC31DOWNTO12_shadow /= EX_ADD_RES32DOWNTO332DOWNTO13_shadow_intermed_1) else '0';
dfp_trap_vector(2759) <= '1' when (V_F_PC31DOWNTO12_shadow /= XC_TRAP_ADDRESS31DOWNTO12_shadow_intermed_1) else '0';
dfp_trap_vector(2760) <= '1' when (V_F_PC31DOWNTO12_shadow /= R.F.PC( 31 DOWNTO 12 )) else '0';
dfp_trap_vector(2761) <= '1' when (V_F_PC31DOWNTO12_shadow /= RIN_M_CTRL_PC31DOWNTO12_intermed_4) else '0';
dfp_trap_vector(2762) <= '1' when (V_F_PC31DOWNTO12_shadow /= IR_ADDR31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(2763) <= '1' when (V_F_PC31DOWNTO12_shadow /= R_X_CTRL_PC31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(2764) <= '1' when (V_F_PC31DOWNTO12_shadow /= R_D_PC31DOWNTO12_intermed_6) else '0';
dfp_trap_vector(2765) <= '1' when (V_F_PC31DOWNTO12_shadow /= RIN_X_CTRL_PC31DOWNTO12_intermed_3) else '0';
dfp_trap_vector(2766) <= '1' when (V_F_PC31DOWNTO12_shadow /= RIN_D_PC31DOWNTO12_intermed_7) else '0';
dfp_trap_vector(2767) <= '1' when (V_F_PC31DOWNTO12_shadow /= VIR_ADDR31DOWNTO12_shadow_intermed_2) else '0';
dfp_trap_vector(2768) <= '1' when (V_F_PC31DOWNTO12_shadow /= V_M_CTRL_PC31DOWNTO12_shadow_intermed_4) else '0';
dfp_trap_vector(2769) <= '1' when (XC_VECTT3DOWNTO0_shadow /= V_X_CTRL_TT3DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(2770) <= '1' when (XC_VECTT3DOWNTO0_shadow /= R_M_CTRL_TT3DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2771) <= '1' when (XC_VECTT3DOWNTO0_shadow /= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(2772) <= '1' when (XC_VECTT3DOWNTO0_shadow /= R_X_RESULT6DOWNTO03DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2773) <= '1' when (XC_VECTT3DOWNTO0_shadow /= R_A_CTRL_TT3DOWNTO0_intermed_3) else '0';
dfp_trap_vector(2774) <= '1' when (XC_VECTT3DOWNTO0_shadow /= RIN_A_CTRL_TT3DOWNTO0_intermed_4) else '0';
dfp_trap_vector(2775) <= '1' when (XC_VECTT3DOWNTO0_shadow /= V_A_CTRL_TT3DOWNTO0_shadow_intermed_4) else '0';
dfp_trap_vector(2776) <= '1' when (XC_VECTT3DOWNTO0_shadow /= R_E_CTRL_TT3DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2777) <= '1' when (XC_VECTT3DOWNTO0_shadow /= RIN_M_CTRL_TT3DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2778) <= '1' when (XC_VECTT3DOWNTO0_shadow /= V_M_CTRL_TT3DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(2779) <= '1' when (XC_VECTT3DOWNTO0_shadow /= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2780) <= '1' when (XC_VECTT3DOWNTO0_shadow /= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2781) <= '1' when (XC_VECTT3DOWNTO0_shadow /= R.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 )) else '0';
dfp_trap_vector(2782) <= '1' when (XC_VECTT3DOWNTO0_shadow /= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(2783) <= '1' when (XC_VECTT3DOWNTO0_shadow /= V_E_CTRL_TT3DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(2784) <= '1' when (XC_VECTT3DOWNTO0_shadow /= RIN_X_CTRL_TT3DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2785) <= '1' when (XC_VECTT3DOWNTO0_shadow /= R.X.CTRL.TT( 3 DOWNTO 0 )) else '0';
dfp_trap_vector(2786) <= '1' when (XC_VECTT3DOWNTO0_shadow /= RIN_E_CTRL_TT3DOWNTO0_intermed_3) else '0';
dfp_trap_vector(2787) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= V_X_CTRL_TT3DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(2788) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= R_M_CTRL_TT3DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2789) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(2790) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= R_X_RESULT6DOWNTO03DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2791) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= R_A_CTRL_TT3DOWNTO0_intermed_4) else '0';
dfp_trap_vector(2792) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= RIN_A_CTRL_TT3DOWNTO0_intermed_5) else '0';
dfp_trap_vector(2793) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= V_A_CTRL_TT3DOWNTO0_shadow_intermed_5) else '0';
dfp_trap_vector(2794) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= R_E_CTRL_TT3DOWNTO0_intermed_3) else '0';
dfp_trap_vector(2795) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= RIN_W_S_TT3DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2796) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= RIN_M_CTRL_TT3DOWNTO0_intermed_3) else '0';
dfp_trap_vector(2797) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= V_M_CTRL_TT3DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(2798) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_3) else '0';
dfp_trap_vector(2799) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2800) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= R.W.S.TT( 3 DOWNTO 0 )) else '0';
dfp_trap_vector(2801) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= R_X_RESULT6DOWNTO03DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2802) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(2803) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= V_E_CTRL_TT3DOWNTO0_shadow_intermed_4) else '0';
dfp_trap_vector(2804) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= RIN_X_CTRL_TT3DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2805) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= R_X_CTRL_TT3DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2806) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= RIN_E_CTRL_TT3DOWNTO0_intermed_4) else '0';
dfp_trap_vector(2807) <= '1' when (V_W_S_TT3DOWNTO0_shadow /= XC_VECTT3DOWNTO0_shadow_intermed_1) else '0';
dfp_trap_vector(2808) <= '1' when (V_A_CTRL_PC31DOWNTO2_shadow /= V_D_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2809) <= '1' when (V_A_CTRL_PC31DOWNTO2_shadow /= RIN_D_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2810) <= '1' when (V_A_CTRL_PC31DOWNTO2_shadow /= R_D_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2811) <= '1' when (V_A_CTRL_PC31DOWNTO2_shadow /= RIN_A_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2812) <= '1' when (V_A_CTRL_PC31DOWNTO2_shadow /= R.A.CTRL.PC( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(2813) <= '1' when (V_X_DATA03_shadow /= V_X_DATA03_shadow_intermed_2) else '0';
dfp_trap_vector(2814) <= '1' when (V_X_DATA03_shadow /= DCO_DATA03_intermed_1) else '0';
dfp_trap_vector(2815) <= '1' when (V_X_DATA03_shadow /= RIN_X_DATA03_intermed_1) else '0';
dfp_trap_vector(2816) <= '1' when (V_X_DATA03_shadow /= R_X_DATA03_intermed_1) else '0';
dfp_trap_vector(2817) <= '1' when (V_X_DATA03_shadow /= RIN_X_DATA03_intermed_2) else '0';
dfp_trap_vector(2818) <= '1' when (V_X_DATA03_shadow /= R.X.DATA ( 0 )( 3 )) else '0';
dfp_trap_vector(2819) <= '1' when (VIR_ADDR31DOWNTO12_shadow /= R_M_CTRL_PC31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(2820) <= '1' when (VIR_ADDR31DOWNTO12_shadow /= V_D_PC31DOWNTO12_shadow_intermed_6) else '0';
dfp_trap_vector(2821) <= '1' when (VIR_ADDR31DOWNTO12_shadow /= V_A_CTRL_PC31DOWNTO12_shadow_intermed_5) else '0';
dfp_trap_vector(2822) <= '1' when (VIR_ADDR31DOWNTO12_shadow /= V_E_CTRL_PC31DOWNTO12_shadow_intermed_4) else '0';
dfp_trap_vector(2823) <= '1' when (VIR_ADDR31DOWNTO12_shadow /= R_A_CTRL_PC31DOWNTO12_intermed_4) else '0';
dfp_trap_vector(2824) <= '1' when (VIR_ADDR31DOWNTO12_shadow /= R_E_CTRL_PC31DOWNTO12_intermed_3) else '0';
dfp_trap_vector(2825) <= '1' when (VIR_ADDR31DOWNTO12_shadow /= RIN_A_CTRL_PC31DOWNTO12_intermed_5) else '0';
dfp_trap_vector(2826) <= '1' when (VIR_ADDR31DOWNTO12_shadow /= RIN_E_CTRL_PC31DOWNTO12_intermed_4) else '0';
dfp_trap_vector(2827) <= '1' when (VIR_ADDR31DOWNTO12_shadow /= IRIN_ADDR31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(2828) <= '1' when (VIR_ADDR31DOWNTO12_shadow /= V_X_CTRL_PC31DOWNTO12_shadow_intermed_2) else '0';
dfp_trap_vector(2829) <= '1' when (VIR_ADDR31DOWNTO12_shadow /= RIN_M_CTRL_PC31DOWNTO12_intermed_3) else '0';
dfp_trap_vector(2830) <= '1' when (VIR_ADDR31DOWNTO12_shadow /= IR.ADDR( 31 DOWNTO 12 )) else '0';
dfp_trap_vector(2831) <= '1' when (VIR_ADDR31DOWNTO12_shadow /= R_X_CTRL_PC31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(2832) <= '1' when (VIR_ADDR31DOWNTO12_shadow /= R_D_PC31DOWNTO12_intermed_5) else '0';
dfp_trap_vector(2833) <= '1' when (VIR_ADDR31DOWNTO12_shadow /= RIN_X_CTRL_PC31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(2834) <= '1' when (VIR_ADDR31DOWNTO12_shadow /= RIN_D_PC31DOWNTO12_intermed_6) else '0';
dfp_trap_vector(2835) <= '1' when (VIR_ADDR31DOWNTO12_shadow /= V_M_CTRL_PC31DOWNTO12_shadow_intermed_3) else '0';
dfp_trap_vector(2836) <= '1' when (VIR_ADDR31DOWNTO2_shadow /= RIN_M_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2837) <= '1' when (VIR_ADDR31DOWNTO2_shadow /= V_D_PC31DOWNTO2_shadow_intermed_6) else '0';
dfp_trap_vector(2838) <= '1' when (VIR_ADDR31DOWNTO2_shadow /= RIN_D_PC31DOWNTO2_intermed_6) else '0';
dfp_trap_vector(2839) <= '1' when (VIR_ADDR31DOWNTO2_shadow /= RIN_X_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2840) <= '1' when (VIR_ADDR31DOWNTO2_shadow /= IRIN_ADDR31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2841) <= '1' when (VIR_ADDR31DOWNTO2_shadow /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(2842) <= '1' when (VIR_ADDR31DOWNTO2_shadow /= R_D_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2843) <= '1' when (VIR_ADDR31DOWNTO2_shadow /= R_M_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2844) <= '1' when (VIR_ADDR31DOWNTO2_shadow /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(2845) <= '1' when (VIR_ADDR31DOWNTO2_shadow /= RIN_A_CTRL_PC31DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2846) <= '1' when (VIR_ADDR31DOWNTO2_shadow /= R_A_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2847) <= '1' when (VIR_ADDR31DOWNTO2_shadow /= V_M_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(2848) <= '1' when (VIR_ADDR31DOWNTO2_shadow /= R_X_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2849) <= '1' when (VIR_ADDR31DOWNTO2_shadow /= R_E_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2850) <= '1' when (VIR_ADDR31DOWNTO2_shadow /= IR.ADDR( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(2851) <= '1' when (VIR_ADDR31DOWNTO2_shadow /= RIN_E_CTRL_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2852) <= '1' when (VIR_ADDR31DOWNTO2_shadow /= V_X_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2853) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= V_F_PC31DOWNTO4_shadow_intermed_1) else '0';
dfp_trap_vector(2854) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= V_X_CTRL_PC31DOWNTO4_shadow_intermed_3) else '0';
dfp_trap_vector(2855) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= IR_ADDR31DOWNTO4_intermed_1) else '0';
dfp_trap_vector(2856) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= R.F.PC( 31 DOWNTO 4 )) else '0';
dfp_trap_vector(2857) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= VIR_ADDR31DOWNTO4_shadow_intermed_2) else '0';
dfp_trap_vector(2858) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= RIN_F_PC31DOWNTO4_intermed_1) else '0';
dfp_trap_vector(2859) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= RIN_A_CTRL_PC31DOWNTO4_intermed_6) else '0';
dfp_trap_vector(2860) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= R_A_CTRL_PC31DOWNTO4_intermed_5) else '0';
dfp_trap_vector(2861) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= R_D_PC31DOWNTO4_intermed_6) else '0';
dfp_trap_vector(2862) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= RIN_X_CTRL_PC31DOWNTO4_intermed_3) else '0';
dfp_trap_vector(2863) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= EX_ADD_RES32DOWNTO332DOWNTO5_shadow_intermed_1) else '0';
dfp_trap_vector(2864) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= V_D_PC31DOWNTO4_shadow_intermed_7) else '0';
dfp_trap_vector(2865) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= V_E_CTRL_PC31DOWNTO4_shadow_intermed_5) else '0';
dfp_trap_vector(2866) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= RIN_M_CTRL_PC31DOWNTO4_intermed_4) else '0';
dfp_trap_vector(2867) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= R_X_CTRL_PC31DOWNTO4_intermed_2) else '0';
dfp_trap_vector(2868) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= IRIN_ADDR31DOWNTO4_intermed_2) else '0';
dfp_trap_vector(2869) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= V_M_CTRL_PC31DOWNTO4_shadow_intermed_4) else '0';
dfp_trap_vector(2870) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= R_M_CTRL_PC31DOWNTO4_intermed_3) else '0';
dfp_trap_vector(2871) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= RIN_D_PC31DOWNTO4_intermed_7) else '0';
dfp_trap_vector(2872) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= RIN_E_CTRL_PC31DOWNTO4_intermed_5) else '0';
dfp_trap_vector(2873) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= EX_JUMP_ADDRESS31DOWNTO4_shadow_intermed_1) else '0';
dfp_trap_vector(2874) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= V_A_CTRL_PC31DOWNTO4_shadow_intermed_6) else '0';
dfp_trap_vector(2875) <= '1' when (XC_TRAP_ADDRESS31DOWNTO4_shadow /= R_E_CTRL_PC31DOWNTO4_intermed_4) else '0';
dfp_trap_vector(2876) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= R_D_PC3DOWNTO2_intermed_6) else '0';
dfp_trap_vector(2877) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= V_D_PC3DOWNTO2_shadow_intermed_7) else '0';
dfp_trap_vector(2878) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= VIR_ADDR3DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2879) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= RIN_D_PC3DOWNTO2_intermed_7) else '0';
dfp_trap_vector(2880) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= R_M_CTRL_PC3DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2881) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= R_E_CTRL_PC3DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2882) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= V_E_CTRL_PC3DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(2883) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= RIN_X_CTRL_PC3DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2884) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= R_A_CTRL_PC3DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2885) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= R.F.PC( 3 DOWNTO 2 )) else '0';
dfp_trap_vector(2886) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= V_X_CTRL_PC3DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(2887) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= RIN_M_CTRL_PC3DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2888) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= IRIN_ADDR3DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2889) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= EX_JUMP_ADDRESS3DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(2890) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= EX_ADD_RES32DOWNTO34DOWNTO3_shadow_intermed_1) else '0';
dfp_trap_vector(2891) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= RIN_A_CTRL_PC3DOWNTO2_intermed_6) else '0';
dfp_trap_vector(2892) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= V_F_PC3DOWNTO2_shadow_intermed_1) else '0';
dfp_trap_vector(2893) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= V_A_CTRL_PC3DOWNTO2_shadow_intermed_6) else '0';
dfp_trap_vector(2894) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= IR_ADDR3DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2895) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= V_M_CTRL_PC3DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(2896) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= R_X_CTRL_PC3DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2897) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= RIN_E_CTRL_PC3DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2898) <= '1' when (XC_TRAP_ADDRESS3DOWNTO2_shadow /= RIN_F_PC3DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2899) <= '1' when (V_M_CTRL_RD7DOWNTO0_shadow /= V_E_CTRL_RD7DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(2900) <= '1' when (V_M_CTRL_RD7DOWNTO0_shadow /= R_E_CTRL_RD7DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2901) <= '1' when (V_M_CTRL_RD7DOWNTO0_shadow /= V_A_CTRL_RD7DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(2902) <= '1' when (V_M_CTRL_RD7DOWNTO0_shadow /= RIN_A_CTRL_RD7DOWNTO0_intermed_3) else '0';
dfp_trap_vector(2903) <= '1' when (V_M_CTRL_RD7DOWNTO0_shadow /= R.M.CTRL.RD ( 7 DOWNTO 0 )) else '0';
dfp_trap_vector(2904) <= '1' when (V_M_CTRL_RD7DOWNTO0_shadow /= R_A_CTRL_RD7DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2905) <= '1' when (V_M_CTRL_RD7DOWNTO0_shadow /= RIN_E_CTRL_RD7DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2906) <= '1' when (V_M_CTRL_RD7DOWNTO0_shadow /= RIN_M_CTRL_RD7DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2907) <= '1' when (V_M_CTRL_PC_shadow /= RIN_D_PC_intermed_4) else '0';
dfp_trap_vector(2908) <= '1' when (V_M_CTRL_PC_shadow /= RIN_A_CTRL_PC_intermed_3) else '0';
dfp_trap_vector(2909) <= '1' when (V_M_CTRL_PC_shadow /= R_A_CTRL_PC_intermed_2) else '0';
dfp_trap_vector(2910) <= '1' when (V_M_CTRL_PC_shadow /= V_E_CTRL_PC_shadow_intermed_2) else '0';
dfp_trap_vector(2911) <= '1' when (V_M_CTRL_PC_shadow /= R.M.CTRL.PC) else '0';
dfp_trap_vector(2912) <= '1' when (V_M_CTRL_PC_shadow /= R_E_CTRL_PC_intermed_1) else '0';
dfp_trap_vector(2913) <= '1' when (V_M_CTRL_PC_shadow /= RIN_M_CTRL_PC_intermed_1) else '0';
dfp_trap_vector(2914) <= '1' when (V_M_CTRL_PC_shadow /= V_A_CTRL_PC_shadow_intermed_3) else '0';
dfp_trap_vector(2915) <= '1' when (V_M_CTRL_PC_shadow /= R_D_PC_intermed_3) else '0';
dfp_trap_vector(2916) <= '1' when (V_M_CTRL_PC_shadow /= RIN_E_CTRL_PC_intermed_2) else '0';
dfp_trap_vector(2917) <= '1' when (V_M_CTRL_PC_shadow /= V_D_PC_shadow_intermed_4) else '0';
dfp_trap_vector(2918) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= RIN_M_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2919) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= V_D_PC31DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(2920) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= RIN_D_PC31DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2921) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(2922) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= R_D_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2923) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= R.M.CTRL.PC( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(2924) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= V_E_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2925) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= RIN_A_CTRL_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2926) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= R_A_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2927) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= R_E_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2928) <= '1' when (V_M_CTRL_PC31DOWNTO2_shadow /= RIN_E_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2929) <= '1' when (V_A_CTRL_INST20_shadow /= RIN_A_CTRL_INST20_intermed_1) else '0';
dfp_trap_vector(2930) <= '1' when (V_A_CTRL_INST20_shadow /= R.A.CTRL.INST ( 20 )) else '0';
dfp_trap_vector(2931) <= '1' when (V_A_CTRL_INST20_shadow /= RIN_A_CTRL_INST20_intermed_2) else '0';
dfp_trap_vector(2932) <= '1' when (V_A_CTRL_INST20_shadow /= V_A_CTRL_INST20_shadow_intermed_2) else '0';
dfp_trap_vector(2933) <= '1' when (V_A_CTRL_INST20_shadow /= DE_INST20_shadow_intermed_1) else '0';
dfp_trap_vector(2934) <= '1' when (V_A_CTRL_INST20_shadow /= R_A_CTRL_INST20_intermed_1) else '0';
dfp_trap_vector(2935) <= '1' when (V_A_CTRL_INST20_shadow /= RIN_A_CTRL_INST20_intermed_1) else '0';
dfp_trap_vector(2936) <= '1' when (V_A_CTRL_INST20_shadow /= DE_INST20_shadow_intermed_1) else '0';
dfp_trap_vector(2937) <= '1' when (V_A_CTRL_INST20_shadow /= R.A.CTRL.INST( 20 )) else '0';
dfp_trap_vector(2938) <= '1' when (V_A_CTRL_INST24_shadow /= R_A_CTRL_INST24_intermed_1) else '0';
dfp_trap_vector(2939) <= '1' when (V_A_CTRL_INST24_shadow /= RIN_A_CTRL_INST24_intermed_2) else '0';
dfp_trap_vector(2940) <= '1' when (V_A_CTRL_INST24_shadow /= R.A.CTRL.INST ( 24 )) else '0';
dfp_trap_vector(2941) <= '1' when (V_A_CTRL_INST24_shadow /= V_A_CTRL_INST24_shadow_intermed_2) else '0';
dfp_trap_vector(2942) <= '1' when (V_A_CTRL_INST24_shadow /= DE_INST24_shadow_intermed_1) else '0';
dfp_trap_vector(2943) <= '1' when (V_A_CTRL_INST24_shadow /= RIN_A_CTRL_INST24_intermed_1) else '0';
dfp_trap_vector(2944) <= '1' when (V_A_CTRL_INST24_shadow /= R.A.CTRL.INST( 24 )) else '0';
dfp_trap_vector(2945) <= '1' when (V_A_CTRL_INST24_shadow /= RIN_A_CTRL_INST24_intermed_1) else '0';
dfp_trap_vector(2946) <= '1' when (V_A_CTRL_INST24_shadow /= DE_INST24_shadow_intermed_1) else '0';
dfp_trap_vector(2947) <= '1' when (V_X_CTRL_PC31DOWNTO4_shadow /= RIN_A_CTRL_PC31DOWNTO4_intermed_4) else '0';
dfp_trap_vector(2948) <= '1' when (V_X_CTRL_PC31DOWNTO4_shadow /= R_A_CTRL_PC31DOWNTO4_intermed_3) else '0';
dfp_trap_vector(2949) <= '1' when (V_X_CTRL_PC31DOWNTO4_shadow /= R_D_PC31DOWNTO4_intermed_4) else '0';
dfp_trap_vector(2950) <= '1' when (V_X_CTRL_PC31DOWNTO4_shadow /= RIN_X_CTRL_PC31DOWNTO4_intermed_1) else '0';
dfp_trap_vector(2951) <= '1' when (V_X_CTRL_PC31DOWNTO4_shadow /= V_D_PC31DOWNTO4_shadow_intermed_5) else '0';
dfp_trap_vector(2952) <= '1' when (V_X_CTRL_PC31DOWNTO4_shadow /= V_E_CTRL_PC31DOWNTO4_shadow_intermed_3) else '0';
dfp_trap_vector(2953) <= '1' when (V_X_CTRL_PC31DOWNTO4_shadow /= RIN_M_CTRL_PC31DOWNTO4_intermed_2) else '0';
dfp_trap_vector(2954) <= '1' when (V_X_CTRL_PC31DOWNTO4_shadow /= R.X.CTRL.PC( 31 DOWNTO 4 )) else '0';
dfp_trap_vector(2955) <= '1' when (V_X_CTRL_PC31DOWNTO4_shadow /= V_M_CTRL_PC31DOWNTO4_shadow_intermed_2) else '0';
dfp_trap_vector(2956) <= '1' when (V_X_CTRL_PC31DOWNTO4_shadow /= R_M_CTRL_PC31DOWNTO4_intermed_1) else '0';
dfp_trap_vector(2957) <= '1' when (V_X_CTRL_PC31DOWNTO4_shadow /= RIN_D_PC31DOWNTO4_intermed_5) else '0';
dfp_trap_vector(2958) <= '1' when (V_X_CTRL_PC31DOWNTO4_shadow /= RIN_E_CTRL_PC31DOWNTO4_intermed_3) else '0';
dfp_trap_vector(2959) <= '1' when (V_X_CTRL_PC31DOWNTO4_shadow /= V_A_CTRL_PC31DOWNTO4_shadow_intermed_4) else '0';
dfp_trap_vector(2960) <= '1' when (V_X_CTRL_PC31DOWNTO4_shadow /= R_E_CTRL_PC31DOWNTO4_intermed_2) else '0';
dfp_trap_vector(2961) <= '1' when (V_X_CTRL_PC3DOWNTO2_shadow /= R_D_PC3DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2962) <= '1' when (V_X_CTRL_PC3DOWNTO2_shadow /= V_D_PC3DOWNTO2_shadow_intermed_5) else '0';
dfp_trap_vector(2963) <= '1' when (V_X_CTRL_PC3DOWNTO2_shadow /= RIN_D_PC3DOWNTO2_intermed_5) else '0';
dfp_trap_vector(2964) <= '1' when (V_X_CTRL_PC3DOWNTO2_shadow /= R_M_CTRL_PC3DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2965) <= '1' when (V_X_CTRL_PC3DOWNTO2_shadow /= R_E_CTRL_PC3DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2966) <= '1' when (V_X_CTRL_PC3DOWNTO2_shadow /= V_E_CTRL_PC3DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(2967) <= '1' when (V_X_CTRL_PC3DOWNTO2_shadow /= RIN_X_CTRL_PC3DOWNTO2_intermed_1) else '0';
dfp_trap_vector(2968) <= '1' when (V_X_CTRL_PC3DOWNTO2_shadow /= R_A_CTRL_PC3DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2969) <= '1' when (V_X_CTRL_PC3DOWNTO2_shadow /= RIN_M_CTRL_PC3DOWNTO2_intermed_2) else '0';
dfp_trap_vector(2970) <= '1' when (V_X_CTRL_PC3DOWNTO2_shadow /= RIN_A_CTRL_PC3DOWNTO2_intermed_4) else '0';
dfp_trap_vector(2971) <= '1' when (V_X_CTRL_PC3DOWNTO2_shadow /= V_A_CTRL_PC3DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(2972) <= '1' when (V_X_CTRL_PC3DOWNTO2_shadow /= V_M_CTRL_PC3DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(2973) <= '1' when (V_X_CTRL_PC3DOWNTO2_shadow /= R.X.CTRL.PC( 3 DOWNTO 2 )) else '0';
dfp_trap_vector(2974) <= '1' when (V_X_CTRL_PC3DOWNTO2_shadow /= RIN_E_CTRL_PC3DOWNTO2_intermed_3) else '0';
dfp_trap_vector(2975) <= '1' when (V_M_CTRL_RD6DOWNTO0_shadow /= RIN_E_CTRL_RD6DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2976) <= '1' when (V_M_CTRL_RD6DOWNTO0_shadow /= RIN_M_CTRL_RD6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2977) <= '1' when (V_M_CTRL_RD6DOWNTO0_shadow /= R_E_CTRL_RD6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2978) <= '1' when (V_M_CTRL_RD6DOWNTO0_shadow /= V_E_CTRL_RD6DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(2979) <= '1' when (V_M_CTRL_RD6DOWNTO0_shadow /= V_A_CTRL_RD6DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(2980) <= '1' when (V_M_CTRL_RD6DOWNTO0_shadow /= R_A_CTRL_RD6DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2981) <= '1' when (V_M_CTRL_RD6DOWNTO0_shadow /= RIN_A_CTRL_RD6DOWNTO0_intermed_3) else '0';
dfp_trap_vector(2982) <= '1' when (V_M_CTRL_RD6DOWNTO0_shadow /= R.M.CTRL.RD( 6 DOWNTO 0 )) else '0';
dfp_trap_vector(2983) <= '1' when (V_E_CTRL_TT_shadow /= RIN_A_CTRL_TT_intermed_2) else '0';
dfp_trap_vector(2984) <= '1' when (V_E_CTRL_TT_shadow /= R_A_CTRL_TT_intermed_1) else '0';
dfp_trap_vector(2985) <= '1' when (V_E_CTRL_TT_shadow /= "000000") else '0';
dfp_trap_vector(2986) <= '1' when (V_E_CTRL_TT_shadow /= R.E.CTRL.TT) else '0';
dfp_trap_vector(2987) <= '1' when (V_E_CTRL_TT_shadow /= RIN_E_CTRL_TT_intermed_1) else '0';
dfp_trap_vector(2988) <= '1' when (V_E_CTRL_TT_shadow /= V_A_CTRL_TT_shadow_intermed_2) else '0';
dfp_trap_vector(2989) <= '1' when (V_X_RESULT6DOWNTO03DOWNTO0_shadow /= V_X_RESULT6DOWNTO03DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(2990) <= '1' when (V_X_RESULT6DOWNTO03DOWNTO0_shadow /= R_X_RESULT6DOWNTO03DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2991) <= '1' when (V_X_RESULT6DOWNTO03DOWNTO0_shadow /= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2992) <= '1' when (V_X_RESULT6DOWNTO03DOWNTO0_shadow /= RIN_X_RESULT6DOWNTO03DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2993) <= '1' when (V_X_RESULT6DOWNTO03DOWNTO0_shadow /= R.X.RESULT ( 6 DOWNTO 0 )( 3 DOWNTO 0 )) else '0';
dfp_trap_vector(2994) <= '1' when (V_X_CTRL_TT3DOWNTO0_shadow /= R_M_CTRL_TT3DOWNTO0_intermed_1) else '0';
dfp_trap_vector(2995) <= '1' when (V_X_CTRL_TT3DOWNTO0_shadow /= R_A_CTRL_TT3DOWNTO0_intermed_3) else '0';
dfp_trap_vector(2996) <= '1' when (V_X_CTRL_TT3DOWNTO0_shadow /= RIN_A_CTRL_TT3DOWNTO0_intermed_4) else '0';
dfp_trap_vector(2997) <= '1' when (V_X_CTRL_TT3DOWNTO0_shadow /= V_A_CTRL_TT3DOWNTO0_shadow_intermed_4) else '0';
dfp_trap_vector(2998) <= '1' when (V_X_CTRL_TT3DOWNTO0_shadow /= R_E_CTRL_TT3DOWNTO0_intermed_2) else '0';
dfp_trap_vector(2999) <= '1' when (V_X_CTRL_TT3DOWNTO0_shadow /= RIN_M_CTRL_TT3DOWNTO0_intermed_2) else '0';
dfp_trap_vector(3000) <= '1' when (V_X_CTRL_TT3DOWNTO0_shadow /= V_M_CTRL_TT3DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(3001) <= '1' when (V_X_CTRL_TT3DOWNTO0_shadow /= V_E_CTRL_TT3DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(3002) <= '1' when (V_X_CTRL_TT3DOWNTO0_shadow /= RIN_X_CTRL_TT3DOWNTO0_intermed_1) else '0';
dfp_trap_vector(3003) <= '1' when (V_X_CTRL_TT3DOWNTO0_shadow /= R.X.CTRL.TT( 3 DOWNTO 0 )) else '0';
dfp_trap_vector(3004) <= '1' when (V_X_CTRL_TT3DOWNTO0_shadow /= RIN_E_CTRL_TT3DOWNTO0_intermed_3) else '0';
dfp_trap_vector(3005) <= '1' when (V_X_CTRL_PC31DOWNTO12_shadow /= R_M_CTRL_PC31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(3006) <= '1' when (V_X_CTRL_PC31DOWNTO12_shadow /= V_D_PC31DOWNTO12_shadow_intermed_5) else '0';
dfp_trap_vector(3007) <= '1' when (V_X_CTRL_PC31DOWNTO12_shadow /= V_A_CTRL_PC31DOWNTO12_shadow_intermed_4) else '0';
dfp_trap_vector(3008) <= '1' when (V_X_CTRL_PC31DOWNTO12_shadow /= V_E_CTRL_PC31DOWNTO12_shadow_intermed_3) else '0';
dfp_trap_vector(3009) <= '1' when (V_X_CTRL_PC31DOWNTO12_shadow /= R_A_CTRL_PC31DOWNTO12_intermed_3) else '0';
dfp_trap_vector(3010) <= '1' when (V_X_CTRL_PC31DOWNTO12_shadow /= R_E_CTRL_PC31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(3011) <= '1' when (V_X_CTRL_PC31DOWNTO12_shadow /= RIN_A_CTRL_PC31DOWNTO12_intermed_4) else '0';
dfp_trap_vector(3012) <= '1' when (V_X_CTRL_PC31DOWNTO12_shadow /= RIN_E_CTRL_PC31DOWNTO12_intermed_3) else '0';
dfp_trap_vector(3013) <= '1' when (V_X_CTRL_PC31DOWNTO12_shadow /= RIN_M_CTRL_PC31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(3014) <= '1' when (V_X_CTRL_PC31DOWNTO12_shadow /= R.X.CTRL.PC( 31 DOWNTO 12 )) else '0';
dfp_trap_vector(3015) <= '1' when (V_X_CTRL_PC31DOWNTO12_shadow /= R_D_PC31DOWNTO12_intermed_4) else '0';
dfp_trap_vector(3016) <= '1' when (V_X_CTRL_PC31DOWNTO12_shadow /= RIN_X_CTRL_PC31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(3017) <= '1' when (V_X_CTRL_PC31DOWNTO12_shadow /= RIN_D_PC31DOWNTO12_intermed_5) else '0';
dfp_trap_vector(3018) <= '1' when (V_X_CTRL_PC31DOWNTO12_shadow /= V_M_CTRL_PC31DOWNTO12_shadow_intermed_2) else '0';
dfp_trap_vector(3019) <= '1' when (V_E_CTRL_RD7DOWNTO0_shadow /= R.E.CTRL.RD ( 7 DOWNTO 0 )) else '0';
dfp_trap_vector(3020) <= '1' when (V_E_CTRL_RD7DOWNTO0_shadow /= V_A_CTRL_RD7DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(3021) <= '1' when (V_E_CTRL_RD7DOWNTO0_shadow /= RIN_A_CTRL_RD7DOWNTO0_intermed_2) else '0';
dfp_trap_vector(3022) <= '1' when (V_E_CTRL_RD7DOWNTO0_shadow /= R_A_CTRL_RD7DOWNTO0_intermed_1) else '0';
dfp_trap_vector(3023) <= '1' when (V_E_CTRL_RD7DOWNTO0_shadow /= RIN_E_CTRL_RD7DOWNTO0_intermed_1) else '0';
dfp_trap_vector(3024) <= '1' when (V_E_CTRL_PC_shadow /= RIN_D_PC_intermed_3) else '0';
dfp_trap_vector(3025) <= '1' when (V_E_CTRL_PC_shadow /= RIN_A_CTRL_PC_intermed_2) else '0';
dfp_trap_vector(3026) <= '1' when (V_E_CTRL_PC_shadow /= R_A_CTRL_PC_intermed_1) else '0';
dfp_trap_vector(3027) <= '1' when (V_E_CTRL_PC_shadow /= R.E.CTRL.PC) else '0';
dfp_trap_vector(3028) <= '1' when (V_E_CTRL_PC_shadow /= V_A_CTRL_PC_shadow_intermed_2) else '0';
dfp_trap_vector(3029) <= '1' when (V_E_CTRL_PC_shadow /= R_D_PC_intermed_2) else '0';
dfp_trap_vector(3030) <= '1' when (V_E_CTRL_PC_shadow /= RIN_E_CTRL_PC_intermed_1) else '0';
dfp_trap_vector(3031) <= '1' when (V_E_CTRL_PC_shadow /= V_D_PC_shadow_intermed_3) else '0';
dfp_trap_vector(3032) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= V_D_PC31DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(3033) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= RIN_D_PC31DOWNTO2_intermed_3) else '0';
dfp_trap_vector(3034) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= V_A_CTRL_PC31DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(3035) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= R_D_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(3036) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= RIN_A_CTRL_PC31DOWNTO2_intermed_2) else '0';
dfp_trap_vector(3037) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= R_A_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(3038) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= R.E.CTRL.PC( 31 DOWNTO 2 )) else '0';
dfp_trap_vector(3039) <= '1' when (V_E_CTRL_PC31DOWNTO2_shadow /= RIN_E_CTRL_PC31DOWNTO2_intermed_1) else '0';
dfp_trap_vector(3040) <= '1' when (V_M_CTRL_PC31DOWNTO4_shadow /= RIN_A_CTRL_PC31DOWNTO4_intermed_3) else '0';
dfp_trap_vector(3041) <= '1' when (V_M_CTRL_PC31DOWNTO4_shadow /= R_A_CTRL_PC31DOWNTO4_intermed_2) else '0';
dfp_trap_vector(3042) <= '1' when (V_M_CTRL_PC31DOWNTO4_shadow /= R_D_PC31DOWNTO4_intermed_3) else '0';
dfp_trap_vector(3043) <= '1' when (V_M_CTRL_PC31DOWNTO4_shadow /= V_D_PC31DOWNTO4_shadow_intermed_4) else '0';
dfp_trap_vector(3044) <= '1' when (V_M_CTRL_PC31DOWNTO4_shadow /= V_E_CTRL_PC31DOWNTO4_shadow_intermed_2) else '0';
dfp_trap_vector(3045) <= '1' when (V_M_CTRL_PC31DOWNTO4_shadow /= RIN_M_CTRL_PC31DOWNTO4_intermed_1) else '0';
dfp_trap_vector(3046) <= '1' when (V_M_CTRL_PC31DOWNTO4_shadow /= R.M.CTRL.PC( 31 DOWNTO 4 )) else '0';
dfp_trap_vector(3047) <= '1' when (V_M_CTRL_PC31DOWNTO4_shadow /= RIN_D_PC31DOWNTO4_intermed_4) else '0';
dfp_trap_vector(3048) <= '1' when (V_M_CTRL_PC31DOWNTO4_shadow /= RIN_E_CTRL_PC31DOWNTO4_intermed_2) else '0';
dfp_trap_vector(3049) <= '1' when (V_M_CTRL_PC31DOWNTO4_shadow /= V_A_CTRL_PC31DOWNTO4_shadow_intermed_3) else '0';
dfp_trap_vector(3050) <= '1' when (V_M_CTRL_PC31DOWNTO4_shadow /= R_E_CTRL_PC31DOWNTO4_intermed_1) else '0';
dfp_trap_vector(3051) <= '1' when (V_M_CTRL_PC3DOWNTO2_shadow /= R_D_PC3DOWNTO2_intermed_3) else '0';
dfp_trap_vector(3052) <= '1' when (V_M_CTRL_PC3DOWNTO2_shadow /= V_D_PC3DOWNTO2_shadow_intermed_4) else '0';
dfp_trap_vector(3053) <= '1' when (V_M_CTRL_PC3DOWNTO2_shadow /= RIN_D_PC3DOWNTO2_intermed_4) else '0';
dfp_trap_vector(3054) <= '1' when (V_M_CTRL_PC3DOWNTO2_shadow /= R.M.CTRL.PC( 3 DOWNTO 2 )) else '0';
dfp_trap_vector(3055) <= '1' when (V_M_CTRL_PC3DOWNTO2_shadow /= R_E_CTRL_PC3DOWNTO2_intermed_1) else '0';
dfp_trap_vector(3056) <= '1' when (V_M_CTRL_PC3DOWNTO2_shadow /= V_E_CTRL_PC3DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(3057) <= '1' when (V_M_CTRL_PC3DOWNTO2_shadow /= R_A_CTRL_PC3DOWNTO2_intermed_2) else '0';
dfp_trap_vector(3058) <= '1' when (V_M_CTRL_PC3DOWNTO2_shadow /= RIN_M_CTRL_PC3DOWNTO2_intermed_1) else '0';
dfp_trap_vector(3059) <= '1' when (V_M_CTRL_PC3DOWNTO2_shadow /= RIN_A_CTRL_PC3DOWNTO2_intermed_3) else '0';
dfp_trap_vector(3060) <= '1' when (V_M_CTRL_PC3DOWNTO2_shadow /= V_A_CTRL_PC3DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(3061) <= '1' when (V_M_CTRL_PC3DOWNTO2_shadow /= RIN_E_CTRL_PC3DOWNTO2_intermed_2) else '0';
dfp_trap_vector(3062) <= '1' when (V_E_CTRL_RD6DOWNTO0_shadow /= RIN_E_CTRL_RD6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(3063) <= '1' when (V_E_CTRL_RD6DOWNTO0_shadow /= R.E.CTRL.RD( 6 DOWNTO 0 )) else '0';
dfp_trap_vector(3064) <= '1' when (V_E_CTRL_RD6DOWNTO0_shadow /= V_A_CTRL_RD6DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(3065) <= '1' when (V_E_CTRL_RD6DOWNTO0_shadow /= R_A_CTRL_RD6DOWNTO0_intermed_1) else '0';
dfp_trap_vector(3066) <= '1' when (V_E_CTRL_RD6DOWNTO0_shadow /= RIN_A_CTRL_RD6DOWNTO0_intermed_2) else '0';
dfp_trap_vector(3067) <= '1' when (V_M_CTRL_TT3DOWNTO0_shadow /= R.M.CTRL.TT( 3 DOWNTO 0 )) else '0';
dfp_trap_vector(3068) <= '1' when (V_M_CTRL_TT3DOWNTO0_shadow /= R_A_CTRL_TT3DOWNTO0_intermed_2) else '0';
dfp_trap_vector(3069) <= '1' when (V_M_CTRL_TT3DOWNTO0_shadow /= RIN_A_CTRL_TT3DOWNTO0_intermed_3) else '0';
dfp_trap_vector(3070) <= '1' when (V_M_CTRL_TT3DOWNTO0_shadow /= V_A_CTRL_TT3DOWNTO0_shadow_intermed_3) else '0';
dfp_trap_vector(3071) <= '1' when (V_M_CTRL_TT3DOWNTO0_shadow /= R_E_CTRL_TT3DOWNTO0_intermed_1) else '0';
dfp_trap_vector(3072) <= '1' when (V_M_CTRL_TT3DOWNTO0_shadow /= RIN_M_CTRL_TT3DOWNTO0_intermed_1) else '0';
dfp_trap_vector(3073) <= '1' when (V_M_CTRL_TT3DOWNTO0_shadow /= V_E_CTRL_TT3DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(3074) <= '1' when (V_M_CTRL_TT3DOWNTO0_shadow /= RIN_E_CTRL_TT3DOWNTO0_intermed_2) else '0';
dfp_trap_vector(3075) <= '1' when (V_M_CTRL_PC31DOWNTO12_shadow /= R.M.CTRL.PC( 31 DOWNTO 12 )) else '0';
dfp_trap_vector(3076) <= '1' when (V_M_CTRL_PC31DOWNTO12_shadow /= V_D_PC31DOWNTO12_shadow_intermed_4) else '0';
dfp_trap_vector(3077) <= '1' when (V_M_CTRL_PC31DOWNTO12_shadow /= V_A_CTRL_PC31DOWNTO12_shadow_intermed_3) else '0';
dfp_trap_vector(3078) <= '1' when (V_M_CTRL_PC31DOWNTO12_shadow /= V_E_CTRL_PC31DOWNTO12_shadow_intermed_2) else '0';
dfp_trap_vector(3079) <= '1' when (V_M_CTRL_PC31DOWNTO12_shadow /= R_A_CTRL_PC31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(3080) <= '1' when (V_M_CTRL_PC31DOWNTO12_shadow /= R_E_CTRL_PC31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(3081) <= '1' when (V_M_CTRL_PC31DOWNTO12_shadow /= RIN_A_CTRL_PC31DOWNTO12_intermed_3) else '0';
dfp_trap_vector(3082) <= '1' when (V_M_CTRL_PC31DOWNTO12_shadow /= RIN_E_CTRL_PC31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(3083) <= '1' when (V_M_CTRL_PC31DOWNTO12_shadow /= RIN_M_CTRL_PC31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(3084) <= '1' when (V_M_CTRL_PC31DOWNTO12_shadow /= R_D_PC31DOWNTO12_intermed_3) else '0';
dfp_trap_vector(3085) <= '1' when (V_M_CTRL_PC31DOWNTO12_shadow /= RIN_D_PC31DOWNTO12_intermed_4) else '0';
dfp_trap_vector(3086) <= '1' when (V_E_CTRL_PC31DOWNTO4_shadow /= RIN_A_CTRL_PC31DOWNTO4_intermed_2) else '0';
dfp_trap_vector(3087) <= '1' when (V_E_CTRL_PC31DOWNTO4_shadow /= R_A_CTRL_PC31DOWNTO4_intermed_1) else '0';
dfp_trap_vector(3088) <= '1' when (V_E_CTRL_PC31DOWNTO4_shadow /= R_D_PC31DOWNTO4_intermed_2) else '0';
dfp_trap_vector(3089) <= '1' when (V_E_CTRL_PC31DOWNTO4_shadow /= V_D_PC31DOWNTO4_shadow_intermed_3) else '0';
dfp_trap_vector(3090) <= '1' when (V_E_CTRL_PC31DOWNTO4_shadow /= RIN_D_PC31DOWNTO4_intermed_3) else '0';
dfp_trap_vector(3091) <= '1' when (V_E_CTRL_PC31DOWNTO4_shadow /= RIN_E_CTRL_PC31DOWNTO4_intermed_1) else '0';
dfp_trap_vector(3092) <= '1' when (V_E_CTRL_PC31DOWNTO4_shadow /= V_A_CTRL_PC31DOWNTO4_shadow_intermed_2) else '0';
dfp_trap_vector(3093) <= '1' when (V_E_CTRL_PC31DOWNTO4_shadow /= R.E.CTRL.PC( 31 DOWNTO 4 )) else '0';
dfp_trap_vector(3094) <= '1' when (V_E_CTRL_PC3DOWNTO2_shadow /= R_D_PC3DOWNTO2_intermed_2) else '0';
dfp_trap_vector(3095) <= '1' when (V_E_CTRL_PC3DOWNTO2_shadow /= V_D_PC3DOWNTO2_shadow_intermed_3) else '0';
dfp_trap_vector(3096) <= '1' when (V_E_CTRL_PC3DOWNTO2_shadow /= RIN_D_PC3DOWNTO2_intermed_3) else '0';
dfp_trap_vector(3097) <= '1' when (V_E_CTRL_PC3DOWNTO2_shadow /= R.E.CTRL.PC( 3 DOWNTO 2 )) else '0';
dfp_trap_vector(3098) <= '1' when (V_E_CTRL_PC3DOWNTO2_shadow /= R_A_CTRL_PC3DOWNTO2_intermed_1) else '0';
dfp_trap_vector(3099) <= '1' when (V_E_CTRL_PC3DOWNTO2_shadow /= RIN_A_CTRL_PC3DOWNTO2_intermed_2) else '0';
dfp_trap_vector(3100) <= '1' when (V_E_CTRL_PC3DOWNTO2_shadow /= V_A_CTRL_PC3DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(3101) <= '1' when (V_E_CTRL_PC3DOWNTO2_shadow /= RIN_E_CTRL_PC3DOWNTO2_intermed_1) else '0';
dfp_trap_vector(3102) <= '1' when (V_E_CTRL_TT3DOWNTO0_shadow /= R_A_CTRL_TT3DOWNTO0_intermed_1) else '0';
dfp_trap_vector(3103) <= '1' when (V_E_CTRL_TT3DOWNTO0_shadow /= RIN_A_CTRL_TT3DOWNTO0_intermed_2) else '0';
dfp_trap_vector(3104) <= '1' when (V_E_CTRL_TT3DOWNTO0_shadow /= V_A_CTRL_TT3DOWNTO0_shadow_intermed_2) else '0';
dfp_trap_vector(3105) <= '1' when (V_E_CTRL_TT3DOWNTO0_shadow /= R.E.CTRL.TT( 3 DOWNTO 0 )) else '0';
dfp_trap_vector(3106) <= '1' when (V_E_CTRL_TT3DOWNTO0_shadow /= RIN_E_CTRL_TT3DOWNTO0_intermed_1) else '0';
dfp_trap_vector(3107) <= '1' when (V_E_CTRL_PC31DOWNTO12_shadow /= V_D_PC31DOWNTO12_shadow_intermed_3) else '0';
dfp_trap_vector(3108) <= '1' when (V_E_CTRL_PC31DOWNTO12_shadow /= V_A_CTRL_PC31DOWNTO12_shadow_intermed_2) else '0';
dfp_trap_vector(3109) <= '1' when (V_E_CTRL_PC31DOWNTO12_shadow /= R_A_CTRL_PC31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(3110) <= '1' when (V_E_CTRL_PC31DOWNTO12_shadow /= R.E.CTRL.PC( 31 DOWNTO 12 )) else '0';
dfp_trap_vector(3111) <= '1' when (V_E_CTRL_PC31DOWNTO12_shadow /= RIN_A_CTRL_PC31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(3112) <= '1' when (V_E_CTRL_PC31DOWNTO12_shadow /= RIN_E_CTRL_PC31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(3113) <= '1' when (V_E_CTRL_PC31DOWNTO12_shadow /= R_D_PC31DOWNTO12_intermed_2) else '0';
dfp_trap_vector(3114) <= '1' when (V_E_CTRL_PC31DOWNTO12_shadow /= RIN_D_PC31DOWNTO12_intermed_3) else '0';
dfp_trap_vector(3115) <= '1' when (V_A_CTRL_PC31DOWNTO4_shadow /= RIN_A_CTRL_PC31DOWNTO4_intermed_1) else '0';
dfp_trap_vector(3116) <= '1' when (V_A_CTRL_PC31DOWNTO4_shadow /= R.A.CTRL.PC( 31 DOWNTO 4 )) else '0';
dfp_trap_vector(3117) <= '1' when (V_A_CTRL_PC31DOWNTO4_shadow /= R_D_PC31DOWNTO4_intermed_1) else '0';
dfp_trap_vector(3118) <= '1' when (V_A_CTRL_PC31DOWNTO4_shadow /= V_D_PC31DOWNTO4_shadow_intermed_2) else '0';
dfp_trap_vector(3119) <= '1' when (V_A_CTRL_PC31DOWNTO4_shadow /= RIN_D_PC31DOWNTO4_intermed_2) else '0';
dfp_trap_vector(3120) <= '1' when (V_A_CTRL_PC3DOWNTO2_shadow /= R_D_PC3DOWNTO2_intermed_1) else '0';
dfp_trap_vector(3121) <= '1' when (V_A_CTRL_PC3DOWNTO2_shadow /= V_D_PC3DOWNTO2_shadow_intermed_2) else '0';
dfp_trap_vector(3122) <= '1' when (V_A_CTRL_PC3DOWNTO2_shadow /= RIN_D_PC3DOWNTO2_intermed_2) else '0';
dfp_trap_vector(3123) <= '1' when (V_A_CTRL_PC3DOWNTO2_shadow /= R.A.CTRL.PC( 3 DOWNTO 2 )) else '0';
dfp_trap_vector(3124) <= '1' when (V_A_CTRL_PC3DOWNTO2_shadow /= RIN_A_CTRL_PC3DOWNTO2_intermed_1) else '0';
dfp_trap_vector(3125) <= '1' when (V_A_CTRL_PC31DOWNTO12_shadow /= V_D_PC31DOWNTO12_shadow_intermed_2) else '0';
dfp_trap_vector(3126) <= '1' when (V_A_CTRL_PC31DOWNTO12_shadow /= R.A.CTRL.PC( 31 DOWNTO 12 )) else '0';
dfp_trap_vector(3127) <= '1' when (V_A_CTRL_PC31DOWNTO12_shadow /= RIN_A_CTRL_PC31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(3128) <= '1' when (V_A_CTRL_PC31DOWNTO12_shadow /= R_D_PC31DOWNTO12_intermed_1) else '0';
dfp_trap_vector(3129) <= '1' when (V_A_CTRL_PC31DOWNTO12_shadow /= RIN_D_PC31DOWNTO12_intermed_2) else '0';

dfp_or_reduce : process(dfp_trap_vector)
	variable or_reduce_1565 : std_logic_vector(1564 downto 0);
	variable or_reduce_783 : std_logic_vector(782 downto 0);
	variable or_reduce_392 : std_logic_vector(391 downto 0);
	variable or_reduce_196 : std_logic_vector(195 downto 0);
	variable or_reduce_98 : std_logic_vector(97 downto 0);
	variable or_reduce_49 : std_logic_vector(48 downto 0);
	variable or_reduce_25 : std_logic_vector(24 downto 0);
	variable or_reduce_13 : std_logic_vector(12 downto 0);
	variable or_reduce_7 : std_logic_vector(6 downto 0);
	variable or_reduce_4 : std_logic_vector(3 downto 0);
	variable or_reduce_2 : std_logic_vector(1 downto 0);
begin
	or_reduce_1565 := dfp_trap_vector(3129 downto 1565) OR dfp_trap_vector(1564 downto 0);
	or_reduce_783 := or_reduce_1565(1564 downto 782) OR ("0" & or_reduce_1565(781 downto 0));
	or_reduce_392 := or_reduce_783(782 downto 391) OR ("0" & or_reduce_783(390 downto 0));
	or_reduce_196 := or_reduce_392(391 downto 196) OR or_reduce_392(195 downto 0);
	or_reduce_98 := or_reduce_196(195 downto 98) OR or_reduce_196(97 downto 0);
	or_reduce_49 := or_reduce_98(97 downto 49) OR or_reduce_98(48 downto 0);
	or_reduce_25 := or_reduce_49(48 downto 24) OR ("0" & or_reduce_49(23 downto 0));
	or_reduce_13 := or_reduce_25(24 downto 12) OR ("0" & or_reduce_25(11 downto 0));
	or_reduce_7 := or_reduce_13(12 downto 6) OR ("0" & or_reduce_13(5 downto 0));
	or_reduce_4 := or_reduce_7(6 downto 3) OR ("0" & or_reduce_7(2 downto 0));
	or_reduce_2 := or_reduce_4(3 downto 2) OR or_reduce_4(1 downto 0);
	or_reduce_1 <= or_reduce_2(0) OR or_reduce_2(1);
end process;

  trap_enable_delay : process(clk)
  begin
    if(rising_edge(clk))then
      if(rstn = '0')then
        dfp_delay_start <= 15;
      elsif(dfp_delay_start /= 0)then
        dfp_delay_start <= dfp_delay_start - 1;
      end if;
    end if;
  end process;

  trap_mem : process(clk)
  begin
    if(rising_edge(clk))then
      if(rstn = '0')then
        dfp_trap_mem <= (others => '0');
      elsif(dfp_delay_start = 0)then
        dfp_trap_mem <= dfp_trap_mem OR dfp_trap_vector;
      end if;
    end if;
  end process;

  handlerTrap <= or_reduce_1 when (dfp_delay_start = 0) else '0';
  preg : process (sclk)
  begin 
    if rising_edge(sclk) then 
      rp <= rpin; 
      if rstn = '0' then rp.error <= '0'; end if;
    end if;
  end process;

  reg : process (clk)
  begin
    if rising_edge(clk) then
      if (holdn = '1') then
        r <= rin;
      else
	r.x.ipend <= rin.x.ipend;
	r.m.werr <= rin.m.werr;
	if (holdn or ico.mds) = '0' then
          r.d.inst <= rin.d.inst; r.d.mexc <= rin.d.mexc; 
          r.d.set <= rin.d.set;
        end if;
	if (holdn or dco.mds) = '0' then
          r.x.data <= rin.x.data; r.x.mexc <= rin.x.mexc; 
          r.x.set <= rin.x.set;
        end if;
      end if;
      if rstn = '0' then
        r.w.s.s <= '1'; r.w.s.ps <= '1'; 
        if need_extra_sync_reset(fabtech) /= 0 then 
          r.d.inst <= (others => (others => '0'));
	  r.x.mexc <= '0';
        end if; 
      end if; 
    end if;
  end process;

    dsureg : process(clk) begin
      if rising_edge(clk) then 
	if holdn = '1' then
          dsur <= dsuin;
        else
          dsur.crdy <= dsuin.crdy;
        end if;
	if holdn = '1' then ir <= irin; end if;
      end if;
    end process;

  dummy <= '1';
end;
